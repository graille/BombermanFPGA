library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.PROJECT_PARAMS_PKG.all;
use work.PROJECT_TYPES_PKG.all;
use work.PROJECT_DIRECTION_PKG.all;

entity characters_sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_id : in block_category_type;
        in_sprite_state : in state_type;
        in_sprite_direction : in direction_type;

        in_sprite_row : in integer range 0 to 39;
        in_sprite_col : in integer range 0 to 39;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end characters_sprite_rom;

architecture behavioral of characters_sprite_rom is
    subtype word_t is std_logic_vector(0 to 199);
    type memory_t is array(0 to 3359) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- 0_character_0_0
                (x"fffffffffffffffffe94a529def7b4a529ffffffffffffffff"),
                (x"fffffffffffffffffe94a529def7b4a529ffffffffffffffff"),
                (x"fffffffffffffffa53ac633ac6319d677b4a5294a7ffffffff"),
                (x"ffffffffffffff4ef58c60d8c18d8cef7ac60d8ced3fffffff"),
                (x"fffffffffffd29d6758318d8318c6ceb18c1b3bda7ffffffff"),
                (x"fffffffffffd28c1b18c60d8318c7d63183677bded3fffffff"),
                (x"fffffffffffd28c1b18c60d8318c7d63183677bded3fffffff"),
                (x"ffffffffffa77ac18d8c60d8c18d8c6318ceb0631b29ffffff"),
                (x"ffffffffffa77bd60d8c6318c18d8c6319d60d8cef7b4a7fff"),
                (x"ffffffffffa77bd6306c6318c6318c6318c677bda529ffffff"),
                (x"ffffffffffa77bd6306c6318c6318c6318c677bda529ffffff"),
                (x"ffffffffffa77bdeb06c6758cef58c6318cef694a529ffffff"),
                (x"ffffffffffa77aceb18c6758cef58ceb18cef7bda529ffffff"),
                (x"ffffffffffa77ac6759def7acef7aceb18ca53bded29ffffff"),
                (x"ffffffffff0528c653bded3acef59da319da5294e83fffffff"),
                (x"ffffffffff0529d677bded3bdef59da77bda7694a03fffffff"),
                (x"ffffffffff0529d677bded3bdef59da77bda7694a03fffffff"),
                (x"fffffffffff8014ef59def7bdef59da529da77bd07ffffffff"),
                (x"fffffffffff8014ed18c6759da53bded294a769407ffffffff"),
                (x"fffffffffffffe0a53ac675c8bdeaeed294a5000ffffffffff"),
                (x"fffffffffffffff0529def50ea51d5ed29da53ffffffffffff"),
                (x"fffffffffffffff0529def50ea51d5ed29da53ffffffffffff"),
                (x"ffffffffffffbcf25294a76b4ef695ed294a11eff7ffffffff"),
                (x"ffffffffff7908109034a75dd633aee80002042123ffffffff"),
                (x"ffffffffff28421094210868c18d940842128421097fffffff"),
                (x"ffffffffef094a523c81093a318c7420424790a5285fffffff"),
                (x"ffffffffef094a523c81093a318c7420424790a5285fffffff"),
                (x"fffffffffe204212bc842069d18fb40908479421093dffffff"),
                (x"ffffffffec4b18cf00a108434633b4084250798c6259ffffff"),
                (x"ffffffffe04dee9053c529094ef684214bee8129ba41ffffff"),
                (x"ffffffffff0000065294a79f4ef5eff5294a3000003fffffff"),
                (x"ffffffffff0000065294a79f4ef5eff5294a3000003fffffff"),
                (x"fffffffffffffff0518c6318ca518c6318ca03ffffffffffff"),
                (x"ffffffffffffffffd18c6318ca518c6318ca7fffffffffffff"),
                (x"ffffffffffffffffd28c63194a528c63194a7fffffffffffff"),
                (x"ffffffffffffffff8294a529400294a529407fffffffffffff"),
                (x"ffffffffffffffff8294a529400294a529407fffffffffffff"),
                (x"ffffffffffffffff8294a3294002946529407fffffffffffff"),
                (x"fffffffffffffffffc0c63180ffc0c63180fffffffffffffff"),
                (x"fffffffffffffffffc1defba0ffc1df77a0fffffffffffffff"),

                -- 0_character_0_1
                (x"fffffffffffffffffe94a53bdef694ed294a7fffffffffffff"),
                (x"fffffffffffffffffe94a53bdef694ed294a7fffffffffffff"),
                (x"fffffffffffffffa53ac63063633bda77bded294ffffffffff"),
                (x"fffffffffffd294eb18318c6318d8cef7b4ef7bda7ffffffff"),
                (x"ffffffffffa77bd6319def58c6306ced29d633bda7ffffffff"),
                (x"fffffffffffd294ed3ac63063633bd677ac60d8ced3fffffff"),
                (x"fffffffffffd294ed3ac63063633bd677ac60d8ced3fffffff"),
                (x"fffffffffffd29def7b4a758318d9da529460c63ed3fffffff"),
                (x"ffffffffffa77bd677bdef68cef5894a534e8d8ced3fffffff"),
                (x"ffffffffffa77acef7ac633b44a537bdee9a0fbded3fffffff"),
                (x"ffffffffffa77acef7ac633b44a537bdee9a0fbded3fffffff"),
                (x"ffffffffffa77aceb06318d89bdef7bdef7a33bda7ffffffff"),
                (x"ffffffffffa77b460d8c677b7bdef7bdef7eb29407ffffffff"),
                (x"ffffffffffa529d677b4a53b7bdd2c63197ef400ffffffffff"),
                (x"ffffffffffa529ded294a77b7bdd2500017ed000ffffffffff"),
                (x"fffffffffffd29da53b7bf7b7bdd2400017a5c00ffffffffff"),
                (x"fffffffffffd29da53b7bf7b7bdd2400017a5c00ffffffffff"),
                (x"fffffffffffd294ef697bf537bdee4ef7b74dc00ffffffffff"),
                (x"ffffffffff739dded294a5137bdee4f7bd7bdc00ffffffffff"),
                (x"ffffffffff72115e8294a5137bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffdeb9c870294a5197bdef7bdef7ba400ffffffffff"),
                (x"fffffffffdeb9c870294a5197bdef7bdef7ba400ffffffffff"),
                (x"ffffffd28c677aea7e94a528cbdef7bdef7483ffffffffffff"),
                (x"ffffffb18ced29ffffc4210be6318c6318007fffffffffffff"),
                (x"ffffffd28ced29fff8810848f295ef6001efffffffffffffff"),
                (x"ffffffd29da7ffff15e52bde5f782163185f7fffffffffffff"),
                (x"ffffffd29da7ffff15e52bde5f782163185f7fffffffffffff"),
                (x"ffffffd29da7ffff3c81084aff7bc165adef7fffffffffffff"),
                (x"ffffffd294ffffff10bef798c0001e2b18cf7fffffffffffff"),
                (x"fffffff7bffffff01597bdd37bdd200daccf7fffffffffffff"),
                (x"fffffffffffffff032f7bdef7bdee025accf7fffffffffffff"),
                (x"fffffffffffffff032f7bdef7bdee025accf7fffffffffffff"),
                (x"ffffffffffffffff8137bdd37bdd202dadefffffffffffffff"),
                (x"fffffffffffffffffc000318c0000c677bffffffffffffffff"),
                (x"fffffffffffffffffc14a5294a518ca77bffffffffffffffff"),
                (x"ffffffffffffffffffe0052946318cefffffffffffffffffff"),
                (x"ffffffffffffffffffe0052946318cefffffffffffffffffff"),
                (x"ffffffffffffffffffe00528c63194ffffffffffffffffffff"),
                (x"fffffffffffffffffffff828c63180ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83be297c0ffffffffffffffffffff"),

                -- 0_character_0_2
                (x"fffffffffffffffffe94a769def594a5294fffffffffffffff"),
                (x"fffffffffffffffffe94a769def594a5294fffffffffffffff"),
                (x"fffffffffffd294a53ac6328c18d9d677bda53ffffffffffff"),
                (x"ffffffffffa77a31b18c633ac18fac1b19def694ffffffffff"),
                (x"fffffffffffd29d60d9def7ac631831b19deb3bda7ffffffff"),
                (x"ffffffffffa77bdeb06c677ac633ac677bd60d8ca7ffffffff"),
                (x"ffffffffffa77bdeb06c677ac633ac677bd60d8ca7ffffffff"),
                (x"fffffffff460c636759def68c18fbded29d18d8ced3fffffff"),
                (x"ffffffd28c1b18c1b3b4a319d18fbda3194eb3bda53fffffff"),
                (x"fffffff7b4a77bd675894dd3d18fbda252cef7bded3fffffff"),
                (x"fffffff7b4a77bd675894dd3d18fbda252cef7bded3fffffff"),
                (x"ffffffd294ed294ed137bdefd18fb462529ef58c653fffffff"),
                (x"fffffffff4ef7bda32f7bdefd633b44dee96518ced3fffffff"),
                (x"fffffffff4eb19da26f7bdefdef689bdef74f7bded3fffffff"),
                (x"ffffffffffa77acedd8c632fda51376318cbd3bda7ffffffff"),
                (x"ffffffffff0529dedca0002f44a6f700005ba694483fffffff"),
                (x"ffffffffff0529dedca0002f44a6f700005ba694483fffffff"),
                (x"ffffffffff025204dc80002e9bdef700004ba400b83fffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"fffffffffffbde5026f7bdef7bdef7bdef7480a57fffffffff"),
                (x"fffffffffffbde5026f7bdef7bdef7bdef7480a57fffffffff"),
                (x"ffffffffff790812b137bdef7bdef7bdee96142123ffffffff"),
                (x"ffffffffef284212158c62537bdee94b18c29021095fffffff"),
                (x"ffffffbde4214af214a10bd8c6318c78425291ef2908f7ffff"),
                (x"fffff794bef1085794a42043ef7bc1090852bca527bc52bfff"),
                (x"fffff794bef1085794a42043ef7bc1090852bca527bc52bfff"),
                (x"fffff7b1894b184f008f785ecb598f0bde4078846252c63fff"),
                (x"fffff62537ba52c000810bca1630a5784240018c4dee94b3ff"),
                (x"fffff625374def7601e10842cb59810842f032f7ba6e94b3ff"),
                (x"ffffff80094def7653cf7908cb598423dfea32f7ba52007fff"),
                (x"ffffff80094def7653cf7908cb598423dfea32f7ba52007fff"),
                (x"ffffffffe04def70519ef7bde633def7bcca02f7ba41ffffff"),
                (x"ffffffffff00000fd18c6318c6318c6318ca7c00003fffffff"),
                (x"fffffffffffffffff68c63194ef68c63194effffffffffffff"),
                (x"ffffffffffffffff828c631940028c6319407fffffffffffff"),
                (x"ffffffffffffffff828c631940028c6319407fffffffffffff"),
                (x"ffffffffffffffff828c631940028c6319407fffffffffffff"),
                (x"fffffffffffffffffc14a5280ffc14a5280fffffffffffffff"),
                (x"ffffffffffffffffffbdefba0ffc1df77bdfffffffffffffff"),

                -- 0_character_0_3
                (x"ffffffffffffffffd29def7bdef7b4a7ffffffffffffffffff"),
                (x"ffffffffffffffffd29def7bdef7b4a7ffffffffffffffffff"),
                (x"fffffa77ac1f7b4a758318d8c6318ced294fffffffffffffff"),
                (x"ffffffd29d60c7d631831b3ac18d9d6319da7fffffffffffff"),
                (x"fffffffff4eb19d6318c675836318c18c63653ffffffffffff"),
                (x"fffffffff4ef7bdeb19deb06c630631b18c67694ffffffffff"),
                (x"fffffffff4ef7bdeb19deb06c630631b18c67694ffffffffff"),
                (x"ffffffd29d6319d60d9def59d63063677bdef694ffffffffff"),
                (x"fffffa77acef7bd1b3b4a33bda53bdeb18c67694ffffffffff"),
                (x"ffffffd29ded28c1b28c6252cef7ac60c631b3bda7ffffffff"),
                (x"ffffffd29ded28c1b28c6252cef7ac60c631b3bda7ffffffff"),
                (x"fffffffff4a52831f5894dee96329deb18c677bda7ffffffff"),
                (x"ffffffffff077a367537bdef74a68c677bd677bda7ffffffff"),
                (x"ffffffffff077acea58c632f7bde9d6319da7694ffffffffff"),
                (x"fffffffffffd29d4dc0001537bdd94a77bded294ffffffffff"),
                (x"fffffffffff8009bdc0001137bdd9ded294ef694ffffffffff"),
                (x"fffffffffff8009bdc0001137bdd9ded294ef694ffffffffff"),
                (x"fffffffffff8017bdfbde92f7bdd34bf7bded000ffffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd34a77b4ef5ce77ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a5280ed50877ffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94a5280721ceef7fffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94a5280721ceef7fffffff"),
                (x"fffffffffffffe04def7bdef763294a001fa3bbd633bffffff"),
                (x"fffffffffffffff0018c6318cf78a427bdfffe94eb29ffffff"),
                (x"fffffffffffffffff80c63de57bc810909effe94eb29ffffff"),
                (x"ffffffffffffffff158c6043e295ef2bde5f7fffa769ffffff"),
                (x"ffffffffffffffff158c6043e295ef2bde5f7fffa769ffffff"),
                (x"ffffffffffffffff7acc607de7bca10908ff7fffff69ffffff"),
                (x"ffffffffffffffff31852f8006319ef14a4f7ffffffbffffff"),
                (x"ffffffffffffffff32c108137bdd37bb18507fffffffffffff"),
                (x"ffffffffffffffff32c4202f7bdef7bdeec07fffffffffffff"),
                (x"ffffffffffffffff32c4202f7bdef7bdeec07fffffffffffff"),
                (x"fffffffffffffffffac528137bdd37ba520fffffffffffffff"),
                (x"ffffffffffffffffffac630006318c0001ffffffffffffffff"),
                (x"ffffffffffffffffffb4a3194a5294a001ffffffffffffffff"),
                (x"fffffffffffffffffffdeb18ca529407ffffffffffffffffff"),
                (x"fffffffffffffffffffdeb18ca529407ffffffffffffffffff"),
                (x"fffffffffffffffffffffd18c6329407ffffffffffffffffff"),
                (x"fffffffffffffffffffff818c63280ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83c5f7ba0ffffffffffffffffffff"),

                -- 0_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a529def7b4a529ffffffffffffffff"),
                (x"fffffffffffffffa53ac633ac6319d677b4a5294a7ffffffff"),
                (x"ffffffffffffff4ef58c60d8c18d8cef7ac60d8ced3fffffff"),
                (x"fffffffffffd29d6758318d8318c6ceb18c1b3bda7ffffffff"),
                (x"fffffffffffd29d6758318d8318c6ceb18c1b3bda7ffffffff"),
                (x"fffffffffffd28c1b18c60d8318c7d63183677bded3fffffff"),
                (x"ffffffffffa77ac18d8c60d8c18d8c6318ceb0631b29ffffff"),
                (x"ffffffffffa77bd60d8c6318c18d8c6319d60d8cef7b4a7fff"),
                (x"ffffffffffa77bd60d8c6318c18d8c6319d60d8cef7b4a7fff"),
                (x"ffffffffffa77bd6306c6318c6318c6318c677bda529ffffff"),
                (x"ffffffffffa77bdeb06c6758cef58c6318cef694a529ffffff"),
                (x"ffffffffffa77aceb18c6758cef58ceb18cef7bda529ffffff"),
                (x"ffffffffffa77ac6759def7acef7aceb18ca53bded29ffffff"),
                (x"ffffffffff0528c653bded3acef59da319da5294e83fffffff"),
                (x"ffffffffff0528c653bded3acef59da319da5294e83fffffff"),
                (x"ffffffffff0529d677bded3bdef59da77bda7694a03fffffff"),
                (x"fffffffffff8014ef59def7bdef59da529da77bd07ffffffff"),
                (x"fffffffffff8014ed18c6759da53bded294a769407ffffffff"),
                (x"fffffffffffffe0a53ac675c8bdeaeed294a5000ffffffffff"),
                (x"fffffffffffffe0a53ac675c8bdeaeed294a5000ffffffffff"),
                (x"ffffffffffffffe0529def50ea51d5ed29da53ffffffffffff"),
                (x"ffffffffffffbc525294a76b4ef695ed294a13deffffffffff"),
                (x"fffffffffff14a421434a75dd6319de800008484f7ffffffff"),
                (x"fffffffffff10852bc210868c18c6c0908508421f7ffffffff"),
                (x"fffffffffff10852bc210868c18c6c0908508421f7ffffffff"),
                (x"fffffffffff14a427824207ac18c6c09085084842fbfffffff"),
                (x"ffffffffff67bdef3c81084346307d0908f2948427bfffffff"),
                (x"ffffffffff0318c03ca420421ef594294af08421f33fffffff"),
                (x"fffffffffff8000079e529484a53b4f7bc0f7bde4b3fffffff"),
                (x"fffffffffff8000079e529484a53b4f7bc0f7bde4b3fffffff"),
                (x"fffffffffffffffff694a3194a5294a529d6252907ffffffff"),
                (x"fffffffffffffffff694a318ca528c6529de8000ffffffffff"),
                (x"fffffffffffffffff7b4a518ca53bdef7a007fffffffffffff"),
                (x"fffffffffffffffffc1ded29463014a001ffffffffffffffff"),
                (x"fffffffffffffffffc1ded29463014a001ffffffffffffffff"),
                (x"ffffffffffffffffffe00758cef40007ffffffffffffffffff"),
                (x"fffffffffffffffffffff83c3f781fffffffffffffffffffff"),
                (x"fffffffffffffffffffff83ddef41fffffffffffffffffffff"),

                -- 0_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a53bdef694ed294a7fffffffffffff"),
                (x"fffffffffffffffa53ac63063633bda77bded294ffffffffff"),
                (x"fffffffffffd294eb18318c6318d8cef7b4ef7bda7ffffffff"),
                (x"ffffffffffa77bd6319def58c6306ced29d633bda7ffffffff"),
                (x"ffffffffffa77bd6319def58c6306ced29d633bda7ffffffff"),
                (x"fffffffffffd294ed3ac63063633bd677ac60d8ced3fffffff"),
                (x"fffffffffffd29def7b4a758318d9da529460c63ed3fffffff"),
                (x"ffffffffffa77bd677bdef68cef5894a534e8d8ced3fffffff"),
                (x"ffffffffffa77bd677bdef68cef5894a534e8d8ced3fffffff"),
                (x"ffffffffffa77acef7ac633b44a537bdee9a0fbded3fffffff"),
                (x"ffffffffffa77aceb06318d89bdef7bdef7a33bda7ffffffff"),
                (x"ffffffffffa77b460d8c677b7bdef7bdef7eb29407ffffffff"),
                (x"ffffffffffa529d677b4a53b7bdd2c63197ef400ffffffffff"),
                (x"ffffffffffa529ded294a77b7bdd2500017ed000ffffffffff"),
                (x"ffffffffffa529ded294a77b7bdd2500017ed000ffffffffff"),
                (x"fffffffffffd29da53b7bf7b7bdd2400017a5c00ffffffffff"),
                (x"fffffffffffd294ef697bf537bdee4ef7b74dc00ffffffffff"),
                (x"ffffffffff739dded294a5137bdee4f7bd7bdc00ffffffffff"),
                (x"ffffffffff72115e8294a5137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffff72115e8294a5137bdef7bdef7bdc00ffffffffff"),
                (x"fffffffff4eb9c870294a5197bdef7bdef7ba400ffffffffff"),
                (x"fffffff7ac677aea7e94a528cbdef7bdef7483ffffffffffff"),
                (x"ffffffd28ced29ff83c5290af6318c6318007fffffffffffff"),
                (x"ffffffd29da7ffff80a420425f79ef7801efffffffffffffff"),
                (x"ffffffd29da7ffff80a420425f79ef7801efffffffffffffff"),
                (x"ffffffd294fffff07884214a47bfc427bcc07fffffffffffff"),
                (x"ffffffd29ffffff078af78421f78be27bcc07fffffffffffff"),
                (x"fffffffffffffff03de4215fef780003de567fffffffffffff"),
                (x"fffffffffffffff03fc52f989632f7b800567fffffffffffff"),
                (x"fffffffffffffff03fc52f989632f7b800567fffffffffffff"),
                (x"fffffffffffffff079e0026f74a6f7b800f67fffffffffffff"),
                (x"fffffffffffffffa03def01374a53765280fffffffffffffff"),
                (x"fffffffffffffffa518c6500c630000529ffffffffffffffff"),
                (x"fffffffffffffff0518c6329400294a7ffffffffffffffffff"),
                (x"fffffffffffffff0518c6329400294a7ffffffffffffffffff"),
                (x"fffffffffffffff0528c652940028c6529ffffffffffffffff"),
                (x"ffffffffffffffff818c6328000014f7bdffffffffffffffff"),
                (x"ffffffffffffffff83bef17c0fffffffffffffffffffffffff"),

                -- 0_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a769def594a5294fffffffffffffff"),
                (x"fffffffffffd294a53ac6328c18d9d677bda53ffffffffffff"),
                (x"ffffffffffa77a31b18c633ac18fac1b19def694ffffffffff"),
                (x"fffffffffffd29d60d9def7ac631831b19deb3bda7ffffffff"),
                (x"fffffffffffd29d60d9def7ac631831b19deb3bda7ffffffff"),
                (x"ffffffffffa77bdeb06c677ac633ac677bd60d8ca7ffffffff"),
                (x"fffffffff460c636759def68c18fbded29d18d8ced3fffffff"),
                (x"ffffffd28c1b18c1b3b4a319d18fbda3194eb3bda53fffffff"),
                (x"ffffffd28c1b18c1b3b4a319d18fbda3194eb3bda53fffffff"),
                (x"fffffff7b4a77bd675894dd3d18fbda252cef7bded3fffffff"),
                (x"ffffffd294ed294ed137bdefd18fb462529ef58c653fffffff"),
                (x"fffffffff4ef7bda32f7bdefd633b44dee96518ced3fffffff"),
                (x"fffffffff4eb19da26f7bdefdef689bdef74f7bded3fffffff"),
                (x"ffffffffffa77acedd8c632fda51376318cbd3bda7ffffffff"),
                (x"ffffffffffa77acedd8c632fda51376318cbd3bda7ffffffff"),
                (x"ffffffffff0529dedca0002f44a6f700005ba694483fffffff"),
                (x"ffffffffff025204dc80002e9bdef700004ba400b83fffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"ffffffffffffbcf026f7bdef7bdef7bdef7483def7ffffffff"),
                (x"ffffffffff794a42b137bdef7bdef7bdee96142127bfffffff"),
                (x"ffffffffef290842158c62537bdee94b18c78484217dffffff"),
                (x"fffffffbc423de5211e10bd8c6318c7908f2bc21090bef7fff"),
                (x"fffffffbc423de5211e10bd8c6318c7908f2bc21090bef7fff"),
                (x"fffffffbcf2908f795e42043ef7bc10908f791ef7bcbef7fff"),
                (x"ffffffb18963de503c8f785ecb598f0bde4781294b3dffffff"),
                (x"ffffffb1894b18c03c810bca1630a578420032f7ba59ffffff"),
                (x"ffffffb197ba520fbca10842cb5981094acbdef74a59ffffff"),
                (x"ffffffb197ba520fbca10842cb5981094acbdef74a59ffffff"),
                (x"ffffffb189bb180fd3def148cb5985f7bccbdd296301ffffff"),
                (x"ffffff80094b19ffd18c6318c6318c652804dd8c003fffffff"),
                (x"ffffffffe00001ffd28c6318ca5294a529400000ffffffffff"),
                (x"fffffffffffffffffe8c6318c63014a5294fffffffffffffff"),
                (x"fffffffffffffffffe8c6318c63014a5294fffffffffffffff"),
                (x"fffffffffffffffffff4a318c6301def7bffffffffffffffff"),
                (x"ffffffffffffffffffe00529def40007ffffffffffffffffff"),
                (x"ffffffffffffffffffffff7beef7ffffffffffffffffffffff"),

                -- 0_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffd29def7bdef7b4a7ffffffffffffffffff"),
                (x"fffffa77ac1f7b4a758318d8c6318ced294fffffffffffffff"),
                (x"ffffffd29d60c7d631831b3ac18d9d6319da7fffffffffffff"),
                (x"fffffffff4eb19d6318c675836318c18c63653ffffffffffff"),
                (x"fffffffff4eb19d6318c675836318c18c63653ffffffffffff"),
                (x"fffffffff4ef7bdeb19deb06c630631b18c67694ffffffffff"),
                (x"ffffffd29d6319d60d9def59d63063677bdef694ffffffffff"),
                (x"fffffa77acef7bd1b3b4a33bda53bdeb18c67694ffffffffff"),
                (x"fffffa77acef7bd1b3b4a33bda53bdeb18c67694ffffffffff"),
                (x"ffffffd29ded28c1b28c6252cef7ac60c631b3bda7ffffffff"),
                (x"fffffffff4a52831f5894dee96329deb18c677bda7ffffffff"),
                (x"ffffffffff077a367537bdef74a68c677bd677bda7ffffffff"),
                (x"ffffffffff077acea58c632f7bde9d6319da7694ffffffffff"),
                (x"fffffffffffd28c4dc0001537bdd94a77bded294ffffffffff"),
                (x"fffffffffffd28c4dc0001537bdd94a77bded294ffffffffff"),
                (x"fffffffffff8009bdc0001137bdd9ded294ef694ffffffffff"),
                (x"fffffffffff8017bdfbde92f7bdd34bf7bded000ffffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd34a77b4ef5ce77ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a5280ed50877ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a5280ed50877ffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94a5280721ceed3fffffff"),
                (x"fffffffffffffe04def7bdef763294a001fa3bbd633bffffff"),
                (x"fffffffffffffff0018c6318c7bca42fbc0ffe94eb29ffffff"),
                (x"fffffffffffffffff80f7bdfe29421214a0fffffa769ffffff"),
                (x"fffffffffffffffff80f7bdfe29421214a0fffffa769ffffff"),
                (x"fffffffffffffff033c4213cf210a52109e07ffffd29ffffff"),
                (x"fffffffffffffff033c4278be08421794be07fffffe9ffffff"),
                (x"fffffffffffffff615e00001ef79e523def07fffffffffffff"),
                (x"fffffffffffffff61417bdeec4a59e2fbcf07fffffffffffff"),
                (x"fffffffffffffff61417bdeec4a59e2fbcf07fffffffffffff"),
                (x"fffffffffffffff63c17bdee9bdee903dfe07fffffffffffff"),
                (x"ffffffffffffffff828c65d29bdd20f7bc0a7fffffffffffff"),
                (x"fffffffffffffffffe800000c6301463194a7fffffffffffff"),
                (x"fffffffffffffffffff4a5280a528c6319407fffffffffffff"),
                (x"fffffffffffffffffff4a5280a528c6319407fffffffffffff"),
                (x"fffffffffffffffffe8c63280a52946529407fffffffffffff"),
                (x"ffffffffffffffffffdef50000028c63180fffffffffffffff"),
                (x"fffffffffffffffffffffffff003c5f77a0fffffffffffffff"),

                -- 0_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a529def7b4a529ffffffffffffffff"),
                (x"fffffffffffffffa53ac633ac6319d677b4a5294a7ffffffff"),
                (x"ffffffffffffff4ef58c60d8c18d8cef7ac60d8ced3fffffff"),
                (x"fffffffffffd29d6758318d8318c6ceb18c1b3bda7ffffffff"),
                (x"fffffffffffd29d6758318d8318c6ceb18c1b3bda7ffffffff"),
                (x"fffffffffffd28c1b18c60d8318c7d63183677bded3fffffff"),
                (x"ffffffffffa77ac18d8c60d8c18d8c6318ceb0631b29ffffff"),
                (x"ffffffffffa77bd60d8c6318c18d8c6319d60d8cef7b4a7fff"),
                (x"ffffffffffa77bd60d8c6318c18d8c6319d60d8cef7b4a7fff"),
                (x"ffffffffffa77bd6306c6318c6318c6318c677bda529ffffff"),
                (x"ffffffffffa77bdeb06c6758cef58c6318cef694a529ffffff"),
                (x"ffffffffffa77aceb18c6758cef58ceb18cef7bda529ffffff"),
                (x"ffffffffffa77ac6759def7acef7aceb18ca53bded29ffffff"),
                (x"ffffffffff0528c653bded3acef59da319da5294e83fffffff"),
                (x"ffffffffff0528c653bded3acef59da319da5294e83fffffff"),
                (x"ffffffffff0529d677bded3bdef59da77bda7694a03fffffff"),
                (x"fffffffffff8014ef59def7bdef59da529da77bd07ffffffff"),
                (x"fffffffffff8014ed18c6759da53bded294a769407ffffffff"),
                (x"fffffffffffffe0a53ac675c8bdeaeed294a5000ffffffffff"),
                (x"fffffffffffffe0a53ac675c8bdeaeed294a5000ffffffffff"),
                (x"fffffffffffffff0529def50ea51d5ed29da53deffffffffff"),
                (x"ffffffffffffffe25294a76b4ef695ed294a10a5f7ffffffff"),
                (x"ffffffffffffbc408494a769d633aee8000290842fbfffffff"),
                (x"ffffffffffffbc1084a4207ac18fb408421794a527bfffffff"),
                (x"ffffffffffffbc1084a4207ac18fb408421794a527bfffffff"),
                (x"fffffffffff14a4084a42058318fb409081f10842fbfffffff"),
                (x"fffffffffff1084295e42058363281084247fbdef33fffffff"),
                (x"ffffffffff67bc1085e5297a3ef681090857818c603fffffff"),
                (x"ffffffffff6253ef781ef7a8ca5084294aff000007ffffffff"),
                (x"ffffffffff6253ef781ef7a8ca5084294aff000007ffffffff"),
                (x"fffffffffff80094b3b4a529da529ded294effffffffffffff"),
                (x"fffffffffffffe0077b4a3194a518c65294effffffffffffff"),
                (x"ffffffffffffffff801def7bda518ca529deffffffffffffff"),
                (x"ffffffffffffffffffe00528063294a77a0fffffffffffffff"),
                (x"ffffffffffffffffffe00528063294a77a0fffffffffffffff"),
                (x"fffffffffffffffffffff8000ef58ce801ffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f787e07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0ef7be07ffffffffffffffffff"),

                -- 0_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a53bdef694ed294a7fffffffffffff"),
                (x"fffffffffffffffa53ac63063633bda77bded294ffffffffff"),
                (x"fffffffffffd294eb18318c6318d8cef7b4ef7bda7ffffffff"),
                (x"ffffffffffa77bd6319def58c6306ced29d633bda7ffffffff"),
                (x"ffffffffffa77bd6319def58c6306ced29d633bda7ffffffff"),
                (x"fffffffffffd294ed3ac63063633bd677ac60d8ced3fffffff"),
                (x"fffffffffffd29def7b4a758318d9da529460c63ed3fffffff"),
                (x"ffffffffffa77bd677bdef68cef5894a534e8d8ced3fffffff"),
                (x"ffffffffffa77bd677bdef68cef5894a534e8d8ced3fffffff"),
                (x"ffffffffffa77acef7ac633b44a537bdee9a0fbded3fffffff"),
                (x"ffffffffffa77aceb06318d89bdef7bdef7a33bda7ffffffff"),
                (x"ffffffffffa77b460d8c677b7bdef7bdef7eb29407ffffffff"),
                (x"ffffffffffa529d677b4a5197bdd2c63197ef400ffffffffff"),
                (x"ffffffffffa529ded294a3197bdd2500017ed000ffffffffff"),
                (x"ffffffffffa529ded294a3197bdd2500017ed000ffffffffff"),
                (x"fffffffffffd29da53b7bb197bdd2400017a5c00ffffffffff"),
                (x"fffffffffffd294ef697bb137bdee4ef7b74dc00ffffffffff"),
                (x"ffffffffff739dded294a5137bdee4f7bd7bdc00ffffffffff"),
                (x"ffffffffff72115ed294a5137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffff72115ed294a5137bdef7bdef7bdc00ffffffffff"),
                (x"fffffffff4eb9c875294a5197bdef7bdef7ba400ffffffffff"),
                (x"fffffffff4677aea5294a528cbdef7bdef7483ffffffffffff"),
                (x"fffffffff4677b4f80a4217de6318c6318007fffffffffffff"),
                (x"fffffffff4ed29f01421091e5211ef4801efffffffffffffff"),
                (x"fffffffff4ed29f01421091e5211ef4801efffffffffffffff"),
                (x"fffffffff4ed29ff3c84204be0842461085f7fffffffffffff"),
                (x"fffffffff4a7fe079021094a57bc2cb7bc567fffffffffffff"),
                (x"fffffffffda7fe02f9ef793cf213cc614be4b3ffffffffffff"),
                (x"ffffffffffa7fe0f26f7ba4002108cb14be483ffffffffffff"),
                (x"ffffffffffa7fe0f26f7ba4002108cb14be483ffffffffffff"),
                (x"fffffffffffffff026f7bdee9f78acb7bc007fffffffffffff"),
                (x"fffffffffffffff03137bdef70018cb5280fffffffffffffff"),
                (x"ffffffffffffffff800c626e90018c6529ffffffffffffffff"),
                (x"ffffffffffffffff8294a0000a5194a529ffffffffffffffff"),
                (x"ffffffffffffffff8294a0000a5194a529ffffffffffffffff"),
                (x"fffffffffffffffff7b4a0000a518c6319ffffffffffffffff"),
                (x"ffffffffffffffff801def4000028cef7a0fffffffffffffff"),
                (x"fffffffffffffffffffffffff003be2fbc0fffffffffffffff"),

                -- 0_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a769def594a5294fffffffffffffff"),
                (x"fffffffffffd294a53ac6328c18d9d677bda53ffffffffffff"),
                (x"ffffffffffa77a31b18c633ac18fac1b19def694ffffffffff"),
                (x"fffffffffffd29d60d9def7ac631831b19deb3bda7ffffffff"),
                (x"fffffffffffd29d60d9def7ac631831b19deb3bda7ffffffff"),
                (x"ffffffffffa77bdeb06c677ac633ac677bd60d8ca7ffffffff"),
                (x"fffffffff460c636759def68c18fbded29d18d8ced3fffffff"),
                (x"ffffffd28c1b18c1b3b4a319d18fbda3194eb3bda53fffffff"),
                (x"ffffffd28c1b18c1b3b4a319d18fbda3194eb3bda53fffffff"),
                (x"fffffff7b4a77bd675894dd3d18fbda252cef7bded3fffffff"),
                (x"ffffffd294ed294ed137bdefd18fb462529ef58c653fffffff"),
                (x"fffffffff4ef7bda32f7bdefd633b44dee96518ced3fffffff"),
                (x"fffffffff4eb19da26f7bdefdef689bdef74f7bded3fffffff"),
                (x"ffffffffffa77acedd8c632fda51376318cbd3bda7ffffffff"),
                (x"ffffffffffa77acedd8c632fda51376318cbd3bda7ffffffff"),
                (x"ffffffffff0529dedca0002f44a6f700005ba694483fffffff"),
                (x"ffffffffff025204dc80002e9bdef700004ba400b83fffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"ffffffffffffbde026f7bdef7bdef7bdef7481eff7ffffffff"),
                (x"fffffffffff10812b137bdef7bdef7bdee9614842bffffffff"),
                (x"fffffffffe290840bd8c62537bdee94b18c29084215fffffff"),
                (x"fffffffbc520421795e423d8c6318c7842f210a57909ef7fff"),
                (x"fffffffbc520421795e423d8c6318c7842f210a57909ef7fff"),
                (x"fffffffbc57bdef23de42043ef7bc10908f2bdef215fef7fff"),
                (x"fffffffffe6252903c8f785ecb598f0bde4780a57b12c67fff"),
                (x"ffffffffec4def7600010bca1630a5784247818c6252c67fff"),
                (x"ffffffffec4a537bdd852842cb5981084257fc004deec67fff"),
                (x"ffffffffec4a537bdd852842cb5981084257fc004deec67fff"),
                (x"ffffffffe063189bdd9ef78acb59842fbdea7c0065d2c67fff"),
                (x"ffffffffff0000cba414a318c6318c6318ca7fff6252007fff"),
                (x"fffffffffffffe000294a5294a518c63194a7fff0001ffffff"),
                (x"fffffffffffffffffe94a52806318c63194fffffffffffffff"),
                (x"fffffffffffffffffe94a52806318c63194fffffffffffffff"),
                (x"fffffffffffffffffffdef7a06318c6529ffffffffffffffff"),
                (x"fffffffffffffffffffff8000ef7b4a001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffef7ddefffffffffffffffffff"),

                -- 0_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffd29def7bdef7b4a7ffffffffffffffffff"),
                (x"fffffa77ac1f7b4a758318d8c6318ced294fffffffffffffff"),
                (x"ffffffd29d60c7d631831b3ac18d9d6319da7fffffffffffff"),
                (x"fffffffff4eb19d6318c675836318c18c63653ffffffffffff"),
                (x"fffffffff4eb19d6318c675836318c18c63653ffffffffffff"),
                (x"fffffffff4ef7bdeb19deb06c630631b18c67694ffffffffff"),
                (x"ffffffd29d6319d60d9def59d63063677bdef694ffffffffff"),
                (x"fffffa77acef7bd1b3b4a33bda53bdeb18c67694ffffffffff"),
                (x"fffffa77acef7bd1b3b4a33bda53bdeb18c67694ffffffffff"),
                (x"ffffffd29ded28c1b28c6252cef7ac60c631b3bda7ffffffff"),
                (x"fffffffff4a52831f5894dee96329deb18c677bda7ffffffff"),
                (x"ffffffffff077a367537bdef74a68c677bd677bda7ffffffff"),
                (x"ffffffffff077acea58c632f7bde9d6319da7694ffffffffff"),
                (x"fffffffffffd29d4dc0001537bdd94a77bded294ffffffffff"),
                (x"fffffffffffd29d4dc0001537bdd94a77bded294ffffffffff"),
                (x"fffffffffff8009bdc0001137bdd9ded294ef694ffffffffff"),
                (x"fffffffffff8017bdfbde92f7bdd34bf7bded000ffffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd34a77b4ef5ce77ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a5280ed50877ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a5280ed50877ffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94a5294721ceefffffffff"),
                (x"fffffffffffffe04def7bdef763294a0014a3bbd677fffffff"),
                (x"fffffffffffffff0018c6318cf7bc5214a0fd3bd653fffffff"),
                (x"fffffffffffffffff8094bde4295e40842507e94ed3fffffff"),
                (x"fffffffffffffffff8094bde4295e40842507e94ed3fffffff"),
                (x"ffffffffffffffff148c61021f78a12108ff7e94ed3fffffff"),
                (x"fffffffffffffff617d6b302f294a508424783ffa53fffffff"),
                (x"fffffffffffffec4f8ac633c47bfc47bdfe283ffff7fffffff"),
                (x"fffffffffffffe04f8b6b308400009bdee9f03ffffffffffff"),
                (x"fffffffffffffe04f8b6b308400009bdee9f03ffffffffffff"),
                (x"fffffffffffffff003d6b30be4a6f7bdee907fffffffffffff"),
                (x"ffffffffffffffff8296b3180bdef7ba52c07fffffffffffff"),
                (x"fffffffffffffffffe8c631804a6e960000fffffffffffffff"),
                (x"fffffffffffffffffe94a519400000a5280fffffffffffffff"),
                (x"fffffffffffffffffe94a519400000a5280fffffffffffffff"),
                (x"fffffffffffffffffd8c6319400000a77bdfffffffffffffff"),
                (x"ffffffffffffffff83bdeb2800001de8000fffffffffffffff"),
                (x"ffffffffffffffff83c52fba0fffffffffffffffffffffffff"),

                -- 1_character_0_0
                (x"fffffffffffffffff7ae739ddef5ce739ddeffffffffffffff"),
                (x"fffffffffffffffff7ae739ddef5ce739ddeffffffffffffff"),
                (x"ffffffffffffffdebab5ad5ce73ab5ad6b573bbdefffffffff"),
                (x"ffffffffffff7aead517ba2aead6b542117456b5777fffffff"),
                (x"ffffffffffffffd73aa84210ead5ceaa108abbbdefffffffff"),
                (x"ffffffffffff7aeadd15ad5ce73ab5756a8ba2b5777fffffff"),
                (x"ffffffffffff7aeadd15ad5ce73ab5756a8ba2b5777fffffff"),
                (x"fffffffffdeb9d5456b5ad6b573915ab9c8ad6b5abbbffffff"),
                (x"fffffff7aead6b5ab9d5aa2b573908ab9d543ab5ad5ddeffff"),
                (x"fffffffffd756b573ab7ba2ae73af7ab9ceaa1ceef7bffffff"),
                (x"fffffffffd756b573ab7ba2ae73af7ab9ceaa1ceef7bffffff"),
                (x"ffffffffffeb9d5abaa8456b5ad6a8756ae756b573bfffffff"),
                (x"fffffffffd756b5756b5ad51573ab5756b573ab5abbbffffff"),
                (x"fffffff7aeab9dd756ae7551573aae739d5739ce739dffffff"),
                (x"fffffef7bdef7ae755ddea2aeef5ceef7ae777bdebbbdeffff"),
                (x"ffffffffff077b573bae722bdef5dd777bd73bbde83fffffff"),
                (x"ffffffffff077b573bae722bdef5dd777bd73bbde83fffffff"),
                (x"ffffffffff077b5777ae755dd73bbd739dd73800e83fffffff"),
                (x"fffffffffff800eebabdebbaead7aeab9dd7740007ffffffff"),
                (x"fffffffffffffe0ebabdef5cead5d5ab9ceef400ffffffffff"),
                (x"fffffffffffffff075ddef5d5739ceab9dde83ffffffffffff"),
                (x"fffffffffffffff075ddef5d5739ceab9dde83ffffffffffff"),
                (x"ffffffffffffffef03ae777aeef7ae739dd07bdeffffffffff"),
                (x"ffffffffffffbc521000077bd003bd70000211eff7ffffffff"),
                (x"fffffffffff14a1084252800000000014a1084212fbfffffff"),
                (x"fffffffffff042109421094a5294a528421284210fbfffffff"),
                (x"fffffffffff042109421094a5294a528421284210fbfffffff"),
                (x"fffffffffe284210f8a1084210842108425f0421097dffffff"),
                (x"fffffffffe294a1280a108421084210842501421297dffffff"),
                (x"fffffffffef14a5078a1084210842108425f00a52fbdffffff"),
                (x"ffffffffff00000f14210842129421084212f800003fffffff"),
                (x"ffffffffff00000f14210842129421084212f800003fffffff"),
                (x"fffffffffffffff0142108421f782108421283ffffffffffff"),
                (x"fffffffffffffffff8a108425f78a10842517fffffffffffff"),
                (x"fffffffffffffffffbdef7bdef7bde1084217fffffffffffff"),
                (x"ffffffffffffffff8047388420004211ce207fffffffffffff"),
                (x"ffffffffffffffff8047388420004211ce207fffffffffffff"),
                (x"ffffffffffffffff804739ce20004739ce207fffffffffffff"),
                (x"fffffffffffffffffc0739ce0ffc0739ce0fffffffffffffff"),
                (x"fffffffffffffffffc14a1280ffc1425280fffffffffffffff"),

                -- 1_character_0_1
                (x"fffffffffffffffffffdef7bdef7bd739ceef7ffffffffffff"),
                (x"fffffffffffffffffffdef7bdef7bd739ceef7ffffffffffff"),
                (x"fffffffffffffffef5ce756b5ad5ce756a8455ce73bfffffff"),
                (x"ffffffffffff7bd756a845ef7422b57210842108abbbffffff"),
                (x"ffffffffffeb9cead508422b5ad6b5ad6b5ab9ceef7fffffff"),
                (x"ffffffffffff7bd756b5ad6f7422ae739d5ad5ceefffffffff"),
                (x"ffffffffffff7bd756b5ad6f7422ae739d5ad5ceefffffffff"),
                (x"ffffffffffeb9cead6a842115739d5ad6ae422b5777fffffff"),
                (x"ffffffffffeb9d5ad508456ae73ab5456bdadef773bbffffff"),
                (x"fffffffffd756b5abab5ab9ce73aa8bb9dd72108ab9ddeffff"),
                (x"fffffffffd756b5abab5ab9ce73aa8bb9dd72108ab9ddeffff"),
                (x"fffffff7aead6ae756ae775ddad508777aced508af7fffffff"),
                (x"fffffffffdeb9ddad5ddeb9dd422aeef7a9ebab5777fffffff"),
                (x"ffffffffffef7b573bae73bb5ad5dd63189676b5efffffffff"),
                (x"ffffffffffeb9ceef7ae775d5739c5000174f5ceefffffffff"),
                (x"ffffffffffef7bdef7bdef5ceef52400017ba7bdffffffffff"),
                (x"ffffffffffef7bdef7bdef5ceef52400017ba7bdffffffffff"),
                (x"ffffffffffef7bdef6894f7a9bdee480017bdc00ffffffffff"),
                (x"ffffffffffff7bdef7b4a5137bdee484217bdc00ffffffffff"),
                (x"ffffffffffff7bdef7bded137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffffffffdf83bded197bdef7bdef7ba400ffffffffff"),
                (x"ffffffffffffffdf83bded197bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffffe9ded28cbdef7bdef7483ffffffffffff"),
                (x"ffffffffffffffffffcf7bde26318c6318007fffffffffffff"),
                (x"fffffffffffffffff8a1084a5297d4a529ffffffffffffffff"),
                (x"fffffffffffffffff82108425084b41dadefffffffffffffff"),
                (x"fffffffffffffffff82108425084b41dadefffffffffffffff"),
                (x"ffffffffffffffff1421094bef78a51b18cfffffffffffffff"),
                (x"ffffffffffffffff04252843e213c5a5296fffffffffffffff"),
                (x"ffffffffffffffff0421084a44a6ec29096fffffffffffffff"),
                (x"fffffffffffffff01421087c34a6ec0d28cfffffffffffffff"),
                (x"fffffffffffffff01421087c34a6ec0d28cfffffffffffffff"),
                (x"ffffffffffffffff80a5297cf63120094befffffffffffffff"),
                (x"fffffffffffffffff80007bde000a1094befffffffffffffff"),
                (x"ffffffffffffffff8bc5294a5084212fbdffffffffffffffff"),
                (x"fffffffffffffffffc4217bdef7bdef7ffffffffffffffffff"),
                (x"fffffffffffffffffc4217bdef7bdef7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0008e739ce0ffffffffffffffffffff"),
                (x"fffffffffffffffffffff804739c40ffffffffffffffffffff"),
                (x"fffffffffffffffffffffd29421280ffffffffffffffffffff"),

                -- 1_character_0_2
                (x"fffffffffffffffff7ae739ceef7ae739ddeffffffffffffff"),
                (x"fffffffffffffffff7ae739ceef7ae739ddeffffffffffffff"),
                (x"ffffffffffff7bd73ab5ad6b5739cead6b5777bdffffffffff"),
                (x"ffffffffffeb9d5aa2e8422b5ad5d545ee8ad5ceefffffffff"),
                (x"ffffffffffff7bd75508455cead5c84211573bbdffffffffff"),
                (x"ffffffffffeb9d545d15abab573bbd756a8bd5ceefffffffff"),
                (x"ffffffffffeb9d545d15abab573bbd756a8bd5ceefffffffff"),
                (x"fffffffffd756b5ad50e756a873baeab9d5aa2b5777bffffff"),
                (x"fffffff7aead6b5722ae7210873bbd456ae756b5ad5ddeffff"),
                (x"fffffffffdef7ae456ae722f773bbd45eee73ab5abbbffffff"),
                (x"fffffffffdef7ae456ae722f773bbd45eee73ab5abbbffffff"),
                (x"ffffffffff739d5abaae755157399d72115eb9ceaf7fffffff"),
                (x"fffffffffd756b5756ae73ab57392ced6b5775ce73bbffffff"),
                (x"ffffffffeeab9ce755ddef5d5ef6e9eb9d5775ce739ddeffff"),
                (x"fffffff7bd777bd73bac633aeef6f7677aeaf5ceef7bdef7ff"),
                (x"ffffffffff077bd774a00013def6f70001d73bbde83fffffff"),
                (x"ffffffffff077bd774a00013def6f70001d73bbde83fffffff"),
                (x"ffffffffff05ee072480002e9ef6f700004eb800b83fffffff"),
                (x"fffffffffff8000edc90802f74a6f7042044f40007ffffffff"),
                (x"fffffffffffffe065c90842f7bdef784204bb000ffffffffff"),
                (x"fffffffffffffff026f7bdef7bdef7bdef7483ffffffffffff"),
                (x"fffffffffffffff026f7bdef7bdef7bdef7483ffffffffffff"),
                (x"fffffffffff7bcff3137bdef7bdef7bdee9679eff7bfffffff"),
                (x"fffffffffe284212f98c62537bdee94b18cf1421097dffffff"),
                (x"fffffffbc5084210fbdef798c6318cf7bdef0421084bef7fff"),
                (x"fffffffbc5294a12f8bef1694632942fbc5f1421294bef7fff"),
                (x"fffffffbc5294a12f8bef1694632942fbc5f1421294bef7fff"),
                (x"ffffff14a10fbc5f78bef04a3b58650fbc5f78a5f04252fbff"),
                (x"ffffff04217908c078252843463281094a1f018c23c210fbff"),
                (x"fffff294a1231974f8210942cb598128421f26f761025297ff"),
                (x"ffffff14a52253749421084a5630a5084212a6f7490a52fbff"),
                (x"ffffff14a52253749421084a5630a5084212a6f7490a52fbff"),
                (x"fffffffbde7b1974942108421294a1084212a6f763fdef7fff"),
                (x"ffffffffff000000142108421f78210842128000003fffffff"),
                (x"ffffffffffffffff80073842100024214a007fffffffffffff"),
                (x"ffffffffffffffff804210842000421084207fffffffffffff"),
                (x"ffffffffffffffff804210842000421084207fffffffffffff"),
                (x"ffffffffffffffff804211c42000423884207fffffffffffff"),
                (x"fffffffffffffffffc0739ce0ffc0739ce0fffffffffffffff"),
                (x"fffffffffffffffffc14a1280ffc1425280fffffffffffffff"),

                -- 1_character_0_3
                (x"ffffffffffffffdeb9ce777bdef7bdefffffffffffffffffff"),
                (x"ffffffffffffffdeb9ce777bdef7bdefffffffffffffffffff"),
                (x"ffffffffee739d5422ae739d5ad6b5739ddeffffffffffffff"),
                (x"fffffff7aeaa1084210e756a8bdef7456b5777bdffffffffff"),
                (x"fffffffffdeb9cead6b5ad6b5ad6a842115ab9ceefffffffff"),
                (x"ffffffffffeb9d5ad5ce73aa8bdef5ad6b5777bdffffffffff"),
                (x"ffffffffffeb9d5ad5ce73aa8bdef5ad6b5777bdffffffffff"),
                (x"fffffffffd756a843ab5ad5cead508456b5ab9ceefffffffff"),
                (x"fffffff7ae75ef7af6a8456ae73ab542115ad5ceefffffffff"),
                (x"fffffeb9ceaa108775d7ba2ae739cead6aead6b5777fffffff"),
                (x"fffffeb9ceaa108775d7ba2ae739cead6aead6b5777fffffff"),
                (x"fffffffffdaa115eb3ae72115ef5dd756b573ab5abbbffffff"),
                (x"fffffffffd756aeea7bdebaa8ef5ceeb9d5af5ceef7fffffff"),
                (x"ffffffffffed6bd6258c675d5ad7ae777ae757bdefffffffff"),
                (x"ffffffffffeb9dd4dc00015cead5dd777bdeb9ceefffffffff"),
                (x"ffffffffffff7a9bdc000113d739ddef7bdef7bdefffffffff"),
                (x"ffffffffffff7a9bdc000113d739ddef7bdef7bdefffffffff"),
                (x"fffffffffff8017bdc10812f74a7bd4d29def7bdefffffffff"),
                (x"fffffffffff8017bde10812f7bdd34a77bdef7bdffffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34ef7bdef7bdffffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94ef7a0ff7ffffffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94ef7a0ff7ffffffffffff"),
                (x"fffffffffffffe04def7bdef763294ed29ffffffffffffffff"),
                (x"fffffffffffffff0018c6318cf79ef7fbdffffffffffffffff"),
                (x"fffffffffffffffffe94a53c5294a1094befffffffffffffff"),
                (x"fffffffffffffffffac31d0a1294210843efffffffffffffff"),
                (x"fffffffffffffffffac31d0a1294210843efffffffffffffff"),
                (x"ffffffffffffffffb183194bef78a508425f7fffffffffffff"),
                (x"ffffffffffffffffda94a17c4f782128421f7fffffffffffff"),
                (x"ffffffffffffffffd8852b2e9210a108421f7fffffffffffff"),
                (x"ffffffffffffffffb1e10b2e918fc10842507fffffffffffff"),
                (x"ffffffffffffffffb1e10b2e918fc10842507fffffffffffff"),
                (x"fffffffffffffffff8a10812c7bfc5294a0fffffffffffffff"),
                (x"fffffffffffffffff8a1084a0f7bde0001efffffffffffffff"),
                (x"ffffffffffffffffffc528421294a52fbdefffffffffffffff"),
                (x"ffffffffffffffffffe210842108421085ffffffffffffffff"),
                (x"ffffffffffffffffffe210842108421085ffffffffffffffff"),
                (x"fffffffffffffffffffff80e739ce207ffffffffffffffffff"),
                (x"fffffffffffffffffffff804739c40ffffffffffffffffffff"),
                (x"fffffffffffffffffffff8284a5280ffffffffffffffffffff"),

                -- 1_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffff7ae739ddef5ce739ddeffffffffffffff"),
                (x"ffffffffffffffdebab5ad5ce73ab5ad6b573bbdefffffffff"),
                (x"ffffffffffff7aead517ba2aead6b542117456b5777fffffff"),
                (x"ffffffffffffffd73aa84210ead5ceaa108abbbdefffffffff"),
                (x"ffffffffffffffd73aa84210ead5ceaa108abbbdefffffffff"),
                (x"ffffffffffff7aeadd15ad5ce73ab5756a8ba2b5777fffffff"),
                (x"fffffffffdeb9d5456b5ad6b573915ab9c8ad6b5abbbffffff"),
                (x"fffffff7aead6b5ab9d5aa2b573908ab9d543ab5ad5ddeffff"),
                (x"fffffff7aead6b5ab9d5aa2b573908ab9d543ab5ad5ddeffff"),
                (x"fffffffffd756b573ab7ba2ae73af7ab9ceaa1ceef7bffffff"),
                (x"ffffffffffeb9d5abaa8456b5ad6a8756ae756b573bfffffff"),
                (x"fffffffffd756b5756b5ad51573ab5756b573ab5abbbffffff"),
                (x"fffffff7aeab9dd756ae7551573aae739d5739ce739dffffff"),
                (x"fffffef7bdef7ae755ddea2aeef5ceef7ae777bdebbbdeffff"),
                (x"fffffef7bdef7ae755ddea2aeef5ceef7ae777bdebbbdeffff"),
                (x"ffffffffff077b573bae722bdef5dd777bd73bbde83fffffff"),
                (x"ffffffffff077b5777ae755dd73bbd739dd73800e83fffffff"),
                (x"fffffffffff800eebabdebbaead7aeab9dd7740007ffffffff"),
                (x"fffffffffffffe0ebabdef5cead5d5ab9ceef400ffffffffff"),
                (x"fffffffffffffe0ebabdef5cead5d5ab9ceef400ffffffffff"),
                (x"fffffffffffffff075ddef5d5739ceab9dde83ffffffffffff"),
                (x"ffffffffffffffe283ae777aeef7ae739dd07bffffffffffff"),
                (x"ffffffffffffbc508400077bd003bd70000097deffffffffff"),
                (x"fffffffffff14a1094252800000000014a1087deffffffffff"),
                (x"fffffffffff14a1094252800000000014a1087deffffffffff"),
                (x"fffffffffff14a52f821094a5294a528425084a5f7ffffffff"),
                (x"ffffffffff294a5f78210842108421094a5084212fbfffffff"),
                (x"ffffffffff014a5f78210842108421094be084212fbfffffff"),
                (x"fffffffffff8000014210842129421094be284212fbfffffff"),
                (x"fffffffffff8000014210842129421094be284212fbfffffff"),
                (x"fffffffffffffff0142108421f78a108425f14a507ffffffff"),
                (x"fffffffffffffff0142108421f78a108425f0000ffffffffff"),
                (x"fffffffffffffff078a5297def7bc5294be07fffffffffffff"),
                (x"fffffffffffffffffc02108e7108421001ffffffffffffffff"),
                (x"fffffffffffffffffc02108e7108421001ffffffffffffffff"),
                (x"ffffffffffffffffffe001e1039c0007ffffffffffffffffff"),
                (x"fffffffffffffffffffff8294a501fffffffffffffffffffff"),
                (x"fffffffffffffffffffff828f18c1fffffffffffffffffffff"),

                -- 1_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffdef7bdef7bd739ceef7ffffffffffff"),
                (x"fffffffffffffffef5ce756b5ad5ce756a8455ce73bfffffff"),
                (x"ffffffffffff7bd756a845ef7422b57210842108abbbffffff"),
                (x"ffffffffffeb9cead508422b5ad6b5ad6b5ab9ceef7fffffff"),
                (x"ffffffffffeb9cead508422b5ad6b5ad6b5ab9ceef7fffffff"),
                (x"ffffffffffff7bd756b5ad6f7422ae739d5ad5ceefffffffff"),
                (x"ffffffffffeb9cead6a842115739d5ad6ae422b5777fffffff"),
                (x"ffffffffffeb9d5ad508456ae73ab5456bdadef773bbffffff"),
                (x"ffffffffffeb9d5ad508456ae73ab5456bdadef773bbffffff"),
                (x"fffffffffd756b5abab5ab9ce73aa8bb9dd72108ab9ddeffff"),
                (x"fffffff7aead6ae756ae775ddad508777aced508af7fffffff"),
                (x"fffffffffdeb9ddad5ddeb9dd422aeef7a9ebab5777fffffff"),
                (x"ffffffffffef7b573bae73bb5ad5dd63189676b5efffffffff"),
                (x"ffffffffffeb9ceef7ae775d5739c5000174f5ceefffffffff"),
                (x"ffffffffffeb9ceef7ae775d5739c5000174f5ceefffffffff"),
                (x"ffffffffffef7bdef7bdef5ceef52400017ba7bdffffffffff"),
                (x"ffffffffffef7bdef6894f7a9bdee480017bdc00ffffffffff"),
                (x"ffffffffffff7bdef7b4a5137bdee484217bdc00ffffffffff"),
                (x"ffffffffffff7bdef7bded137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffffff7bdef7bded137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffffffffdf83bded197bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffffe9ded28cbdef7bdef7483ffffffffffff"),
                (x"ffffffffffffffffffdef14a26318c6318007fffffffffffff"),
                (x"ffffffffffffffffffc528425f7bde1001ffffffffffffffff"),
                (x"ffffffffffffffffffc528425f7bde1001ffffffffffffffff"),
                (x"ffffffffffffffff80a108425294a1a1080fffffffffffffff"),
                (x"ffffffffffffffff80a10842518fde10c6cfffffffffffffff"),
                (x"fffffffffffffff078a1084a121189b842cfffffffffffffff"),
                (x"fffffffffffffff017c52842121197b800cfffffffffffffff"),
                (x"fffffffffffffff017c52842121197b800cfffffffffffffff"),
                (x"ffffffffffffffff17c5294a118d89b8002fffffffffffffff"),
                (x"fffffffffffffff294bef78a52946c00842fffffffffffffff"),
                (x"ffffffffffffffff78a52fbdef780010840fffffffffffffff"),
                (x"ffffffffffffffff7800078a5297de1001ffffffffffffffff"),
                (x"ffffffffffffffff7800078a5297de1001ffffffffffffffff"),
                (x"fffffffffffffff008f081c42000021085ffffffffffffffff"),
                (x"ffffffffffffffff80f0840e0ffc14a529ffffffffffffffff"),
                (x"ffffffffffffffffd294a5080fffffffffffffffffffffffff"),

                -- 1_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffff7ae739ceef7ae739ddeffffffffffffff"),
                (x"ffffffffffff7bd73ab5ad6b5739cead6b5777bdffffffffff"),
                (x"ffffffffffeb9d5aa2e8422b5ad5d545ee8ad5ceefffffffff"),
                (x"ffffffffffff7bd75508455cead5c84211573bbdffffffffff"),
                (x"ffffffffffff7bd75508455cead5c84211573bbdffffffffff"),
                (x"ffffffffffeb9d545d15abab573bbd756a8bd5ceefffffffff"),
                (x"fffffffffd756b5ad50e756a873baeab9d5aa2b5777bffffff"),
                (x"fffffff7aead6b5722ae7210873bbd456ae756b5ad5ddeffff"),
                (x"fffffff7aead6b5722ae7210873bbd456ae756b5ad5ddeffff"),
                (x"fffffffffdef7ae456ae722f773bbd45eee73ab5abbbffffff"),
                (x"ffffffffff739d5abaae755157399d72115eb9ceaf7fffffff"),
                (x"fffffffffd756b5756ae73ab57392ced6b5775ce73bbffffff"),
                (x"ffffffffeeab9ce755ddef5d5ef6e9eb9d5775ce739ddeffff"),
                (x"fffffff7bd777bd73bac633aeef6f7677aeaf5ceef7bdef7ff"),
                (x"fffffff7bd777bd73bac633aeef6f7677aeaf5ceef7bdef7ff"),
                (x"ffffffffff077bd774a00013def6f70001d73bbde83fffffff"),
                (x"ffffffffff05ee072480002e9ef6f700004eb800b83fffffff"),
                (x"fffffffffff8000edc90802f74a6f7042044f40007ffffffff"),
                (x"fffffffffffffe065c90842f7bdef784204bb000ffffffffff"),
                (x"fffffffffffffe065c90842f7bdef784204bb000ffffffffff"),
                (x"fffffffffffffff026f7bdef7bdef7bdef7483ffffffffffff"),
                (x"ffffffffffffbc5f3137bdef7bdef7bdee9678a5f7ffffffff"),
                (x"ffffffffff284212f98c62537bdee94b18c284212fbfffffff"),
                (x"fffffffffe28421094bef798c6318cf7bde08421097dffffff"),
                (x"fffffffffe28421094bef798c6318cf7bde08421097dffffff"),
                (x"fffffffbc5294a12f8252969463294294a5094a5097dffffff"),
                (x"fffffffbc5294a5f14a1084a3b5865094be28421297dffffff"),
                (x"ffffff94a5294be014a5284b4632850842320421097dffffff"),
                (x"fffffffbc420c6000421094acb59852b197490a50fbfffffff"),
                (x"fffffffbc420c6000421094acb59852b197490a50fbfffffff"),
                (x"ffffffbde34bde0f042108421630a10b197b8ca5283fffffff"),
                (x"ffffff800c4b19ff142108421294a1094a948ca507ffffffff"),
                (x"ffffffffe00001fff8a5297de003c52fbde00000ffffffffff"),
                (x"ffffffffffffffff8002108e739c421084207fffffffffffff"),
                (x"ffffffffffffffff8002108e739c421084207fffffffffffff"),
                (x"fffffffffffffffffc0211e1039c4210000fffffffffffffff"),
                (x"ffffffffffffffffffe0040e21080007ffffffffffffffffff"),
                (x"fffffffffffffffffffff82942101fffffffffffffffffffff"),

                -- 1_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffdeb9ce777bdef7bdefffffffffffffffffff"),
                (x"ffffffffee739d5422ae739d5ad6b5739ddeffffffffffffff"),
                (x"fffffff7aeaa1084210e756a8bdef7456b5777bdffffffffff"),
                (x"fffffffffdeb9cead6b5ad6b5ad6a842115ab9ceefffffffff"),
                (x"fffffffffdeb9cead6b5ad6b5ad6a842115ab9ceefffffffff"),
                (x"ffffffffffeb9d5ad5ce73aa8bdef5ad6b5777bdffffffffff"),
                (x"fffffffffd756a843ab5ad5cead508456b5ab9ceefffffffff"),
                (x"fffffff7ae75ef7af6a8456ae73ab542115ad5ceefffffffff"),
                (x"fffffff7ae75ef7af6a8456ae73ab542115ad5ceefffffffff"),
                (x"fffffeb9ceaa108775d7ba2ae739cead6aead6b5777fffffff"),
                (x"fffffffffdaa115eb3ae72115ef5dd756b573ab5abbbffffff"),
                (x"fffffffffd756aeea7bdebaa8ef5ceeb9d5af5ceef7fffffff"),
                (x"ffffffffffed6bd6258c675d5ad7ae777ae757bdefffffffff"),
                (x"ffffffffffeb9dd4dc00015cead5dd777bdeb9ceefffffffff"),
                (x"ffffffffffeb9dd4dc00015cead5dd777bdeb9ceefffffffff"),
                (x"ffffffffffff7a9bdc000113d739ddef7bdef7bdefffffffff"),
                (x"fffffffffff8017bdc10812f74a7bd4d29def7bdefffffffff"),
                (x"fffffffffff8017bde10812f7bdd34a77bdef7bdffffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34ef7bdef7bdffffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34ef7bdef7bdffffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94ef7a0ff7ffffffffffff"),
                (x"fffffffffffffe04def7bdef763294ed29ffffffffffffffff"),
                (x"fffffffffffffff0018c6318cf78a51085ffffffffffffffff"),
                (x"fffffffffffffffffc1ef7bde294212fbdffffffffffffffff"),
                (x"fffffffffffffffffc1ef7bde294212fbdffffffffffffffff"),
                (x"ffffffffffffffff8094a04a529421094a0fffffffffffffff"),
                (x"ffffffffffffffffb07ef7bc329421094a0fffffffffffffff"),
                (x"ffffffffffffffffb037ba584084a1094be07fffffffffffff"),
                (x"ffffffffffffffffb017bdd84084212fbc507fffffffffffff"),
                (x"ffffffffffffffffb017bdd84084212fbc507fffffffffffff"),
                (x"fffffffffffffffff817ba583084a52fbc5f7fffffffffffff"),
                (x"fffffffffffffffffbc003065294bef14a52ffffffffffffff"),
                (x"ffffffffffffffff83def001ef7bde294bef7fffffffffffff"),
                (x"fffffffffffffffffc0217bc5294be0001ef7fffffffffffff"),
                (x"fffffffffffffffffc0217bc5294be0001ef7fffffffffffff"),
                (x"fffffffffffffffffc42108001084781ce207fffffffffffff"),
                (x"fffffffffffffffffe94a501f000f081ce0fffffffffffffff"),
                (x"fffffffffffffffffffffffff00094a5280fffffffffffffff"),

                -- 1_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffff7ae739ddef5ce739ddeffffffffffffff"),
                (x"ffffffffffffffdebab5ad5ce73ab5ad6b573bbdefffffffff"),
                (x"ffffffffffff7aead517ba2aead6b542117456b5777fffffff"),
                (x"ffffffffffffffd73aa84210ead5ceaa108abbbdefffffffff"),
                (x"ffffffffffffffd73aa84210ead5ceaa108abbbdefffffffff"),
                (x"ffffffffffff7aeadd15ad5ce73ab5756a8ba2b5777fffffff"),
                (x"fffffffffdeb9d5456b5ad6b573915ab9c8ad6b5abbbffffff"),
                (x"fffffff7aead6b5ab9d5aa2b573908ab9d543ab5ad5ddeffff"),
                (x"fffffff7aead6b5ab9d5aa2b573908ab9d543ab5ad5ddeffff"),
                (x"fffffffffd756b573ab7ba2ae73af7ab9ceaa1ceef7bffffff"),
                (x"ffffffffffeb9d5abaa8456b5ad6a8756ae756b573bfffffff"),
                (x"fffffffffd756b5756b5ad51573ab5756b573ab5abbbffffff"),
                (x"fffffff7aeab9dd756ae7551573aae739d5739ce739dffffff"),
                (x"fffffef7bdef7ae755ddea2aeef5ceef7ae777bdebbbdeffff"),
                (x"fffffef7bdef7ae755ddea2aeef5ceef7ae777bdebbbdeffff"),
                (x"ffffffffff077b573bae722bdef5dd777bd73bbde83fffffff"),
                (x"ffffffffff077b5777ae755dd73bbd739dd73800e83fffffff"),
                (x"fffffffffff800eebabdebbaead7aeab9dd7740007ffffffff"),
                (x"fffffffffffffe0ebabdef5cead5d5ab9ceef400ffffffffff"),
                (x"fffffffffffffe0ebabdef5cead5d5ab9ceef400ffffffffff"),
                (x"fffffffffffffff075ddef5d5739ceab9dde83ffffffffffff"),
                (x"fffffffffffffff103ae777aeef7ae739dd017deffffffffff"),
                (x"ffffffffffffffe28400077bd003bd70000084a5f7ffffffff"),
                (x"ffffffffffffffe084252800000000014a1284212fbfffffff"),
                (x"ffffffffffffffe084252800000000014a1284212fbfffffff"),
                (x"ffffffffffffbc5084a1094a5294a528421f14a52fbfffffff"),
                (x"fffffffffff14a1084a5284210842108421f78a5297fffffff"),
                (x"fffffffffff14a1087c5284210842108421f78a5283fffffff"),
                (x"fffffffffff14a1097c52842129421084212800007ffffffff"),
                (x"fffffffffff14a1097c52842129421084212800007ffffffff"),
                (x"fffffffffff80052f8a108425f782108421283ffffffffffff"),
                (x"fffffffffffffe0078a108425f782108421283ffffffffffff"),
                (x"ffffffffffffffff83c5294bef7bde294a5103ffffffffffff"),
                (x"ffffffffffffffffffe000842108e710840fffffffffffffff"),
                (x"ffffffffffffffffffe000842108e710840fffffffffffffff"),
                (x"fffffffffffffffffffff800039e103801ffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a529407ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe018df407ffffffffffffffffff"),

                -- 1_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffdef7bdef7bd739ceef7ffffffffffff"),
                (x"fffffffffffffffef5ce756b5ad5ce756a8455ce73bfffffff"),
                (x"ffffffffffff7bd756a845ef7422b57210842108abbbffffff"),
                (x"ffffffffffeb9cead508422b5ad6b5ad6b5ab9ceef7fffffff"),
                (x"ffffffffffeb9cead508422b5ad6b5ad6b5ab9ceef7fffffff"),
                (x"ffffffffffff7bd756b5ad6f7422ae739d5ad5ceefffffffff"),
                (x"ffffffffffeb9cead6a842115739d5ad6ae422b5777fffffff"),
                (x"ffffffffffeb9d5ad508456ae73ab5456bdadef773bbffffff"),
                (x"ffffffffffeb9d5ad508456ae73ab5456bdadef773bbffffff"),
                (x"fffffffffd756b5abab5ab9ce73aa8bb9dd72108ab9ddeffff"),
                (x"fffffff7aead6ae756ae775ddad508777aced508af7fffffff"),
                (x"fffffffffdeb9ddad5ddeb9dd422aeef7a9ebab5777fffffff"),
                (x"ffffffffffef7b573bae73bb5ad5dd63189676b5efffffffff"),
                (x"ffffffffffeb9ceef7ae775d5739c5000174f5ceefffffffff"),
                (x"ffffffffffeb9ceef7ae775d5739c5000174f5ceefffffffff"),
                (x"ffffffffffef7bdef7bdef5ceef52400017ba7bdffffffffff"),
                (x"ffffffffffef7bdef6894f7a9bdee480017bdc00ffffffffff"),
                (x"ffffffffffff7bdef7b4a5137bdee484217bdc00ffffffffff"),
                (x"ffffffffffff7bdef7bded137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffffff7bdef7bded137bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffffffffdf83bded197bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffffe9ded28cbdef7bdef7483ffffffffffff"),
                (x"ffffffffffffffff83c5297de6318c6318007fffffffffffff"),
                (x"fffffffffffffff078a108425f7bd4a529ffffffffffffffff"),
                (x"fffffffffffffff078a108425f7bd4a529ffffffffffffffff"),
                (x"ffffffffffffffff142109421f7823b0c74fffffffffffffff"),
                (x"fffffffffffffe0284252f8a1f78346319467fffffffffffff"),
                (x"fffffffffffffe0284a1087c529425a5ade4b3ffffffffffff"),
                (x"fffffffffffffe02942108483f78a12319e483ffffffffffff"),
                (x"fffffffffffffe02942108483f78a12319e483ffffffffffff"),
                (x"fffffffffffffff014a109077633c5a14be07fffffffffffff"),
                (x"fffffffffffffff078a529197633c1094befffffffffffffff"),
                (x"fffffffffffffff1000210d89000a12fbdefffffffffffffff"),
                (x"fffffffffffffff1084210802108421085ffffffffffffffff"),
                (x"fffffffffffffff1084210802108421085ffffffffffffffff"),
                (x"ffffffffffffffff884000000108e73885ffffffffffffffff"),
                (x"ffffffffffffffff8294a53e01084213de0fffffffffffffff"),
                (x"fffffffffffffffffffffffffa5294a1080fffffffffffffff"),

                -- 1_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffff7ae739ceef7ae739ddeffffffffffffff"),
                (x"ffffffffffff7bd73ab5ad6b5739cead6b5777bdffffffffff"),
                (x"ffffffffffeb9d5aa2e8422b5ad5d545ee8ad5ceefffffffff"),
                (x"ffffffffffff7bd75508455cead5c84211573bbdffffffffff"),
                (x"ffffffffffff7bd75508455cead5c84211573bbdffffffffff"),
                (x"ffffffffffeb9d545d15abab573bbd756a8bd5ceefffffffff"),
                (x"fffffffffd756b5ad50e756a873baeab9d5aa2b5777bffffff"),
                (x"fffffff7aead6b5722ae7210873bbd456ae756b5ad5ddeffff"),
                (x"fffffff7aead6b5722ae7210873bbd456ae756b5ad5ddeffff"),
                (x"fffffffffdef7ae456ae722f773bbd45eee73ab5abbbffffff"),
                (x"ffffffffff739d5abaae755157399d72115eb9ceaf7fffffff"),
                (x"fffffffffd756b5756ae73ab57392ced6b5775ce73bbffffff"),
                (x"ffffffffeeab9ce755ddef5d5ef6e9eb9d5775ce739ddeffff"),
                (x"fffffff7bd777bd73bac633aeef6f7677aeaf5ceef7bdef7ff"),
                (x"fffffff7bd777bd73bac633aeef6f7677aeaf5ceef7bdef7ff"),
                (x"ffffffffff077bd774a00013def6f70001d73bbde83fffffff"),
                (x"ffffffffff05ee072480002e9ef6f700004eb800b83fffffff"),
                (x"fffffffffff8000edc90802f74a6f7042044f40007ffffffff"),
                (x"fffffffffffffe065c90842f7bdef784204bb000ffffffffff"),
                (x"fffffffffffffe065c90842f7bdef784204bb000ffffffffff"),
                (x"fffffffffffffff026f7bdef7bdef7bdef7483ffffffffffff"),
                (x"ffffffffffffbc5f3137bdef7bdef7bdee9678a5f7ffffffff"),
                (x"fffffffffff14a10958c62537bdee94b18cf1421097fffffff"),
                (x"fffffffffe28421087def798c6318cf7bc528421097dffffff"),
                (x"fffffffffe28421087def798c6318cf7bc528421097dffffff"),
                (x"fffffffffe28425284a52969463294294a1f1421294bef7fff"),
                (x"fffffffffe294a1097c5284a3b5865084252f8a5294bef7fff"),
                (x"fffffffffe2842109061084b463285094a5283de294a52ffff"),
                (x"fffffffffff0425226ec614acb598528421080001909ef7fff"),
                (x"fffffffffff0425226ec614acb598528421080001909ef7fff"),
                (x"ffffffffff014a51deec6042563021084210f8007a46f7ffff"),
                (x"fffffffffff80051a5252842529421084212fbff6258007fff"),
                (x"fffffffffffffe0003def14be003de294a5f7fff0001ffffff"),
                (x"ffffffffffffffff80421084239ce71084007fffffffffffff"),
                (x"ffffffffffffffff80421084239ce71084007fffffffffffff"),
                (x"fffffffffffffffffc000084239e1038840fffffffffffffff"),
                (x"fffffffffffffffffffff8000108478001ffffffffffffffff"),
                (x"ffffffffffffffffffffffff42129407ffffffffffffffffff"),

                -- 1_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffdeb9ce777bdef7bdefffffffffffffffffff"),
                (x"ffffffffee739d5422ae739d5ad6b5739ddeffffffffffffff"),
                (x"fffffff7aeaa1084210e756a8bdef7456b5777bdffffffffff"),
                (x"fffffffffdeb9cead6b5ad6b5ad6a842115ab9ceefffffffff"),
                (x"fffffffffdeb9cead6b5ad6b5ad6a842115ab9ceefffffffff"),
                (x"ffffffffffeb9d5ad5ce73aa8bdef5ad6b5777bdffffffffff"),
                (x"fffffffffd756a843ab5ad5cead508456b5ab9ceefffffffff"),
                (x"fffffff7ae75ef7af6a8456ae73ab542115ad5ceefffffffff"),
                (x"fffffff7ae75ef7af6a8456ae73ab542115ad5ceefffffffff"),
                (x"fffffeb9ceaa108775d7ba2ae739cead6aead6b5777fffffff"),
                (x"fffffffffdaa115eb3ae72115ef5dd756b573ab5abbbffffff"),
                (x"fffffffffd756aeea7bdebaa8ef5ceeb9d5af5ceef7fffffff"),
                (x"ffffffffffed6bd6258c675d5ad7ae777ae757bdefffffffff"),
                (x"ffffffffffeb9dd4dc00015cead5dd777bdeb9ceefffffffff"),
                (x"ffffffffffeb9dd4dc00015cead5dd777bdeb9ceefffffffff"),
                (x"ffffffffffff7a9bdc000113d739ddef7bdef7bdefffffffff"),
                (x"fffffffffff8017bdc10812f74a7bd4d29def7bdefffffffff"),
                (x"fffffffffff8017bde10812f7bdd34a77bdef7bdffffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34ef7bdef7bdffffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34ef7bdef7bdffffffffff"),
                (x"fffffffffff8009bdef7bdef7bdd94ef7a0ff7ffffffffffff"),
                (x"fffffffffffffe04def7bdef763294ed29ffffffffffffffff"),
                (x"fffffffffffffff0018c6318cf7bc73fbc0fffffffffffffff"),
                (x"fffffffffffffffffe94a53de29421094be07fffffffffffff"),
                (x"fffffffffffffffffe94a53de29421094be07fffffffffffff"),
                (x"ffffffffffffffffd076b0c3e0842508425f7fffffffffffff"),
                (x"fffffffffffffff6518c6503e084be28421283ffffffffffff"),
                (x"fffffffffffffec4fad4a1425297c1094a1283ffffffffffff"),
                (x"fffffffffffffe04f984204be18c8108425283ffffffffffff"),
                (x"fffffffffffffe04f984204be18c8108425283ffffffffffff"),
                (x"fffffffffffffff078af797ccbdc64094a507fffffffffffff"),
                (x"fffffffffffffffff8a1087ccbdd84294be07fffffffffffff"),
                (x"fffffffffffffffffbc5284a04a583f000017fffffffffffff"),
                (x"fffffffffffffffffc4210842108021084217fffffffffffff"),
                (x"fffffffffffffffffc4210842108021084217fffffffffffff"),
                (x"fffffffffffffffffc4739ce20000000842fffffffffffffff"),
                (x"ffffffffffffffff81e210842003f4a5280fffffffffffffff"),
                (x"ffffffffffffffff8094a5280fffffffffffffffffffffffff"),

                -- 2_character_0_0
                (x"ffffffffffffffffffee739ce739ce739dffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce739dffffffffffffffff"),
                (x"ffffffffffffffffd6b5ad6b573ab5756b577fffffffffffff"),
                (x"fffffffffffffeead517bd6a8ad515aa108ad5ceffffffffff"),
                (x"fffffffffffb9d5422a845eb74211542115aa2b577ffffffff"),
                (x"fffffffffffd6a8ba115add17422a8456a842108afffffffff"),
                (x"fffffffffffd6a8ba115add17422a8456a842108afffffffff"),
                (x"ffffffffff72117ba10842108422a842108422f7abbfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d08abbfffffff"),
                (x"fffffffffdadef7422f7bdd17bdd17bdef7ba108ad7bffffff"),
                (x"fffffffffdadef7422f7bdd17bdd17bdef7ba108ad7bffffff"),
                (x"fffffffffd45ee84210845ef7bdef7bdee842108ad7bffffff"),
                (x"ffffffffee42108421084211742108ba115422b5455dffffff"),
                (x"fffffff7b54210842108421084210842115422b5456bdeffff"),
                (x"fffffff7a8456a8422a8421084210842115422b543abdeffff"),
                (x"ffffffb9c8456a8422a8421084210842115422b543aae77fff"),
                (x"ffffffb9c8456a8422a8421084210842115422b543aae77fff"),
                (x"ffffffb9c8456a8aa2a8422a8ad5084211545508abaae77fff"),
                (x"fffffff7b5439c8aa2b5aa2a8ad508456ae45508ababdeffff"),
                (x"fffffff7ae439d5aa2b5aa2a8ad508456ae43908755ddeffff"),
                (x"fffffffffdaf7b5722ae722a8ad6a8ab9d5abab5757bffffff"),
                (x"fffffffffdaf7b5722ae722a8ad6a8ab9d5abab5757bffffff"),
                (x"ffffffffff077bd756ae755d573ab5777b573bbde83fffffff"),
                (x"ffffffffffffff4ef5cc63baeef5ddeb19def694ffffffffff"),
                (x"fffffffffffd2852b1c42118c6318c2108e6118ca7ffffffff"),
                (x"ffffffffffa14a425084210842108421084a10842d3fffffff"),
                (x"ffffffffffa14a425084210842108421084a10842d3fffffff"),
                (x"ffffffffff714a42d0a4210210842121085a14842bbfffffff"),
                (x"fffffffff4094a528284210842108421094014a52869ffffff"),
                (x"ffffffd28e28424702852908421084214b403884095d4a7fff"),
                (x"ffffffd284094a507ca4210210842121085f80a528494a7fff"),
                (x"ffffffd284094a507ca4210210842121085f80a528494a7fff"),
                (x"ffffffffe07042400084210210842121084000840b81ffffff"),
                (x"ffffffffe04a520fd1c421021084212108ea7c004a41ffffff"),
                (x"ffffffffff0001ffd3bef7bdef7bdef7bdda7fff003fffffff"),
                (x"ffffffffffffffffd3bdefbdef7bdef77bda7fffffffffffff"),
                (x"ffffffffffffffffd3bdefbdef7bdef77bda7fffffffffffff"),
                (x"ffffffffffffffff819defbac0019df77ac07fffffffffffff"),
                (x"fffffffffffffffffc1de8fa0ffc1d1f7a0fffffffffffffff"),
                (x"fffffffffffffffffc0c65980ffc0cb3180fffffffffffffff"),

                -- 2_character_0_1
                (x"fffffffffffffffffdce739d5ad6b5739cefffffffffffffff"),
                (x"fffffffffffffffffdce739d5ad6b5739cefffffffffffffff"),
                (x"fffffffffffffff73aa8422f7bdd15aa11573bffffffffffff"),
                (x"fffffffffffffeeaa117bdef7bdef7ba10845eb5ffffffffff"),
                (x"fffffffffffb9d545508422b5ad6a8bdee8aa2f777ffffffff"),
                (x"ffffffffff756a8aa115ad508bdd15aa117456f7afffffffff"),
                (x"ffffffffff756a8aa115ad508bdd15aa117456f7afffffffff"),
                (x"ffffffffff756b5422a842117422a94b9d5ad5ceabbfffffff"),
                (x"ffffffffeead6b54550845508ad537bdee973929abbfffffff"),
                (x"ffffffffeead6a842115ad6e8ad6f7bdef7bdd29abbfffffff"),
                (x"ffffffffeead6a842115ad6e8ad6f7bdef7bdd29abbfffffff"),
                (x"ffffffffeead6a8aa115aa2f54a6f7bdef7bdd2977ffffffff"),
                (x"ffffffb9d5ab9c8aa2b5aa2f5bdef7bdef7bdd8cefffffffff"),
                (x"ffffffb9d5ab9c8722ae72115bdd2c63197bdc00ffffffffff"),
                (x"ffffffb9d5756a8722ae75515bdd2500017bdc00ffffffffff"),
                (x"fffffff7b5756b5755d7bd50ebdd2400017bdc00ffffffffff"),
                (x"fffffff7b5756b5755d7bd50ebdd2400017bdc00ffffffffff"),
                (x"fffffff7b5756b5757a94b90ebdee439cf7bdc00ffffffffff"),
                (x"fffffff7aeeb9d5757b4a3aaebdee491cf7bdc00ffffffffff"),
                (x"fffffffffda77ae757bdeb9c9bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffffd29d73bbded1c9bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffd29d73bbded1c9bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffa7694a528c4a6f7bdef7483ffffffffffff"),
                (x"fffffffffffffffffe94a168e6318c6318007fffffffffffff"),
                (x"fffffffffffffffffe8420484a50b4a1094a13ffffffffffff"),
                (x"ffffffffffffffffd0a420494210850b9d4f53ffffffffffff"),
                (x"ffffffffffffffffd0a420494210850b9d4f53ffffffffffff"),
                (x"ffffffffffffffffd0a421094a5021239d4f53ffffffffffff"),
                (x"ffffffffffffffffd0a4210b42948109094f7fffffffffffff"),
                (x"fffffffffffffffa3a85294942948429094f53ffffffffffff"),
                (x"fffffffffffffffa1481084852948128434f53ffffffffffff"),
                (x"fffffffffffffffa1481084852948128434f53ffffffffffff"),
                (x"fffffffffffffffa38a529085210212043df53ffffffffffff"),
                (x"ffffffffffffffffd02109004084840f7bdf53ffffffffffff"),
                (x"ffffffffffffffffd1894dc1def421f7bdd07fffffffffffff"),
                (x"fffffffffffffffffc00003bdef7deef7a0fffffffffffffff"),
                (x"fffffffffffffffffc00003bdef7deef7a0fffffffffffffff"),
                (x"ffffffffffffffffffe00018c631800001ffffffffffffffff"),
                (x"fffffffffffffffffffff819ef7ba0ffffffffffffffffffff"),
                (x"fffffffffffffffffffff818cb5980ffffffffffffffffffff"),

                -- 2_character_0_2
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"ffffffffffffffffd6b5ad6b573ab5ad6ae77fffffffffffff"),
                (x"fffffffffffffeead6a845ef5ad517ba108ab9ceffffffffff"),
                (x"fffffffffffb9d545ef7ba117422f7bdef7422b577ffffffff"),
                (x"fffffffffffd6a84210845ee8422f7456b542108afffffffff"),
                (x"fffffffffffd6a84210845ee8422f7456b542108afffffffff"),
                (x"ffffffffff756b545ef7ba11742115aa117ba108abbfffffff"),
                (x"ffffffffff756b5ad6a845dd5422a8bdee8456b5abbfffffff"),
                (x"fffffffffdad6a8455c94dd2ead5c9ba52eaa2b5ad7bffffff"),
                (x"fffffffffdad6a8455c94dd2ead5c9ba52eaa2b5ad7bffffff"),
                (x"fffffffffdaa108bb937bdef7bdef7bdee972108ad7bffffff"),
                (x"ffffffffee456b7abaf7bdef7bdef7bdef775508755dffffff"),
                (x"fffffff7aeab9d7abaf7bdef7bdef7bdef7756f7755ddeffff"),
                (x"fffffff7aeaf7a87258c632f7bdef76318c4baf7ebabdeffff"),
                (x"fffffff7b57252875ca0002f7bdef700005bb9084babdeffff"),
                (x"fffffff7b57252875ca0002f7bdef700005bb9084babdeffff"),
                (x"fffffff7b575ef575c80002f7bdef700004bbab5bbabdeffff"),
                (x"fffffff7b5e8015edc8739ef7bdef739ce4bf6b5075ddeffff"),
                (x"fffffff7aee800e05c9291ef7bdef73ca44b81ce075ddeffff"),
                (x"fffffff7aee801d026f7bdef7bdef7bdef7483bd075ddeffff"),
                (x"fffffff7aee801d026f7bdef7bdef7bdef7483bd075ddeffff"),
                (x"fffffffffd07fe003137bdef7bdef7bdee960000f83bffffff"),
                (x"ffffffffffffff42d00c62537bdee94b180a3294ffffffffff"),
                (x"fffffffffffd285215c52b18c6318c614ae290a5a7ffffffff"),
                (x"ffffffffffa14a4250842109ef7bc421084a10842d3fffffff"),
                (x"ffffffffffa14a4250842109ef7bc421084a10842d3fffffff"),
                (x"ffffffffff714a42d0a10843ef7bc108425a14842bbfffffff"),
                (x"fffffffff4094a5280a42043ef7bc109085014a52869ffffff"),
                (x"ffffffd28e28424702852909ef7bc4214b403884095d4a7fff"),
                (x"ffffffd284094a507ca42109ef7bc421085f80a528494a7fff"),
                (x"ffffffd284094a507ca42109ef7bc421085f80a528494a7fff"),
                (x"ffffffffe070424000842043ef7bc109084000840b81ffffff"),
                (x"ffffffffe04a520fd08108434ef68108424a7c004a41ffffff"),
                (x"ffffffffff0001ffd3a42069def7b40909da7fff003fffffff"),
                (x"ffffffffffffffffd3bdefbddef7bef77bda7fffffffffffff"),
                (x"ffffffffffffffffd3bdefbddef7bef77bda7fffffffffffff"),
                (x"ffffffffffffffff819ef7bac0019df7bcc07fffffffffffff"),
                (x"fffffffffffffffffc1de8fa0ffc1d1f7a0fffffffffffffff"),
                (x"fffffffffffffffffc0c65980ffc0cb3180fffffffffffffff"),

                -- 2_character_0_3
                (x"ffffffffffffffffb9ce756b5ad5ce739dffffffffffffffff"),
                (x"ffffffffffffffffb9ce756b5ad5ce739dffffffffffffffff"),
                (x"fffffffffffffee75515ad517bdee8456ae77fffffffffffff"),
                (x"fffffffffffd6b742117bdef7bdef7ba108abbffffffffffff"),
                (x"ffffffffff75ee8aa2f7ba2b5ad6a842115455ceffffffffff"),
                (x"ffffffffffadef545d15ad51742115aa108aa2b577ffffffff"),
                (x"ffffffffffadef545d15ad51742115aa108aa2b577ffffffff"),
                (x"ffffffffeeab9d5ad5c94a6a8bdd08456a8456b577ffffffff"),
                (x"ffffffffeeaa52e726f7bdd354211542115456b5abbfffffff"),
                (x"ffffffffeeaa537bdef7bdef5422f5aa108422b5abbfffffff"),
                (x"ffffffffeeaa537bdef7bdef5422f5aa108422b5abbfffffff"),
                (x"ffffffffff72537bdef7bdee9ad6e8aa108aa2b5abbfffffff"),
                (x"ffffffffffeb197bdef7bdef7ad6e8ad6a8aa1cead5dffffff"),
                (x"fffffffffff8017bdd8c63137ad508756a8721cead5dffffff"),
                (x"fffffffffff8017bdc0001537ad515756a8722b5755dffffff"),
                (x"fffffffffff8017bdc000113773915bb9d5756b5757bffffff"),
                (x"fffffffffff8017bdc000113773915bb9d5756b5757bffffff"),
                (x"fffffffffff8017bdce7392f77390e4f7b5756b5757bffffff"),
                (x"fffffffffff8017bdcf2912f773aaea77b5755ceebbbffffff"),
                (x"fffffffffff8017bdef7bdef74a5ceef7b573bbda77fffffff"),
                (x"fffffffffff8009bdef7bdef74a5d4ef7ae77694ffffffffff"),
                (x"fffffffffff8009bdef7bdef74a5d4ef7ae77694ffffffffff"),
                (x"fffffffffffffe04def7bdee963294a529da7fffffffffffff"),
                (x"fffffffffffffff0018c6318c73a8ca529ffffffffffffffff"),
                (x"fffffffffffffe4a5094a50b4210812529ffffffffffffffff"),
                (x"ffffffffffffff4f51c109484a5081214b4fffffffffffffff"),
                (x"ffffffffffffff4f51c109484a5081214b4fffffffffffffff"),
                (x"ffffffffffffff4f51c420434a5084214b4fffffffffffffff"),
                (x"ffffffffffffffff508108485a50a4214b4fffffffffffffff"),
                (x"ffffffffffffff4f508529085a50852d28ea7fffffffffffff"),
                (x"ffffffffffffff4f5025284852948109085a7fffffffffffff"),
                (x"ffffffffffffff4f5025284852948109085a7fffffffffffff"),
                (x"ffffffffffffff4f74242042429484294aea7fffffffffffff"),
                (x"ffffffffffffff4f77a1090812100408434fffffffffffffff"),
                (x"fffffffffffffff077def043def4174b194fffffffffffffff"),
                (x"ffffffffffffffff83bdefbddef7a00001ffffffffffffffff"),
                (x"ffffffffffffffff83bdefbddef7a00001ffffffffffffffff"),
                (x"fffffffffffffffffc000018c6318007ffffffffffffffffff"),
                (x"fffffffffffffffffffff83bef7980ffffffffffffffffffff"),
                (x"fffffffffffffffffffff819663180ffffffffffffffffffff"),

                -- 2_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce739dffffffffffffffff"),
                (x"ffffffffffffffffd6b5ad6b573ab5756b577fffffffffffff"),
                (x"fffffffffffffeead517bd6a8ad515aa108ad5ceffffffffff"),
                (x"fffffffffffb9d5422a845eb74211542115aa2b577ffffffff"),
                (x"fffffffffffb9d5422a845eb74211542115aa2b577ffffffff"),
                (x"fffffffffffd6a8ba115add17422a8456a842108afffffffff"),
                (x"ffffffffff72117ba10842108422a842108422f7abbfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d08abbfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d08abbfffffff"),
                (x"fffffffffdadef7422f7bdd17bdd17bdef7ba108ad7bffffff"),
                (x"fffffffffd45ee84210845ef7bdef7bdee842108ad5dffffff"),
                (x"ffffffffee42108421084211742108ba108422b5456bdeffff"),
                (x"fffffff7ae4210842108421084210842115422b543aae77fff"),
                (x"fffffff7b54210842108421084210842115422b543ab5affff"),
                (x"fffffff7b54210842108421084210842115422b543ab5affff"),
                (x"ffffffb9d5456a842108421084210842115421ce455d5abbff"),
                (x"ffffffb9d5456a842115aa108422a84210eaa1ceaa1d5af7ff"),
                (x"ffffffffee4211545515aa115422a84210eaa1ce721ce777ff"),
                (x"fffffffffdaa10e45515ad515422b54210e755ce755ddeffff"),
                (x"fffffffffdaa10e45515ad515422b54210e755ce755ddeffff"),
                (x"ffffffffffed6aead515ab915422ae456ae755ceef41ffffff"),
                (x"ffffffffffff7bdebab5abaaead6bdab9dd73bbdffffffffff"),
                (x"ffffffffffffff423bae715dd739ddef7a5ef694ffffffffff"),
                (x"fffffffffffd284215c42108421084214a5210a5ffffffffff"),
                (x"fffffffffffd284215c42108421084214a5210a5ffffffffff"),
                (x"ffffffffffa10852d0a420421084247528421084a7ffffffff"),
                (x"ffffffffee214a4750a4214a5294a42d2852048477ffffffff"),
                (x"ffffffffe071085a00a421084210842d28e210a5a53fffffff"),
                (x"ffffffffe04b18e0508108421084212528021421203fffffff"),
                (x"ffffffffe04b18e0508108421084212528021421203fffffff"),
                (x"ffffffffff03180038810842121021214ae2058c603fffffff"),
                (x"ffffffffffffffffb88427bde21024739dd03129603fffffff"),
                (x"ffffffffffffffff83def318c003bdef7a0f800007ffffffff"),
                (x"fffffffffffffffffc1de8c7d0000c6001ffffffffffffffff"),
                (x"fffffffffffffffffc1de8c7d0000c6001ffffffffffffffff"),
                (x"ffffffffffffffffffec677cc0000c6001ffffffffffffffff"),
                (x"fffffffffffffffffd8c65acc0000007ffffffffffffffffff"),
                (x"fffffffffffffffffc0c6318c003ffffffffffffffffffffff"),

                -- 2_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffdce739d5ad6b5739cefffffffffffffff"),
                (x"fffffffffffffff73aa8422f7bdd15aa11573bffffffffffff"),
                (x"fffffffffffffeeaa117bdef7bdef7ba10845eb5ffffffffff"),
                (x"fffffffffffb9d545508422b5ad6a8bdee8aa2f777ffffffff"),
                (x"fffffffffffb9d545508422b5ad6a8bdee8aa2f777ffffffff"),
                (x"ffffffffff756a8aa115ad508bdd15aa117456f7afffffffff"),
                (x"ffffffffff756b5422a842117422a94b9d5ad5ceabbfffffff"),
                (x"ffffffffeead6a84550845508ad537bdee973929abbfffffff"),
                (x"ffffffffeead6a84550845508ad537bdee973929abbfffffff"),
                (x"ffffffffeeaa108aa115ad6e8ad6f7bdef7bdd29abbfffffff"),
                (x"ffffffb9d5aa115aa2ae722f54a6f7bdef7bdd2977ffffffff"),
                (x"ffffffb9d5456ae455ce722f5bdef7bdef7bdd8cefffffffff"),
                (x"fffffed6b5456ae455ce72115bdd2c63197bdc00ffffffffff"),
                (x"fffffed6aeab9d5ab9ce75515bdd2500017bdc00ffffffffff"),
                (x"fffffed6aeab9d5ab9ce75515bdd2500017bdc00ffffffffff"),
                (x"fffffed6aeab9d5775d7bd50ebdd2400017bdc00ffffffffff"),
                (x"fffffff7ae739d5ef7a94b90ebdee439cf7bdc00ffffffffff"),
                (x"fffffff7aeeb9d5ebbb4a3aaebdee491cf7bdc00ffffffffff"),
                (x"fffffffffda77aeebbbdeb9c9bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffda77aeebbbdeb9c9bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffffd29debbbded1c9bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffa7694a528c4a6f7bdef7483ffffffffffff"),
                (x"fffffffffffffffffe94a14b46318c6318007fffffffffffff"),
                (x"fffffffffffffffffe8529024210842fbd4fffffffffffffff"),
                (x"fffffffffffffffffe8529024210842fbd4fffffffffffffff"),
                (x"ffffffffffffffffd0a529021294810fbd4fffffffffffffff"),
                (x"ffffffffffffffffd0a529081210a52fbdea7fffffffffffff"),
                (x"ffffffffffffffffd0ae71485210a427bdea7fffffffffffff"),
                (x"fffffffffffffffa14b4a1021210a40fbdea7fffffffffffff"),
                (x"fffffffffffffffa14b4a1021210a40fbdea7fffffffffffff"),
                (x"fffffffffffffff714b4a5081085c40fbdea7fffffffffffff"),
                (x"fffffffffffffffeb894a1021a52810fbdea7fffffffffffff"),
                (x"fffffffffffffffef7a423a89bde840f7bdfffffffffffffff"),
                (x"fffffffffffffff0758c675ce2109def7bdfffffffffffffff"),
                (x"fffffffffffffff0758c675ce2109def7bdfffffffffffffff"),
                (x"fffffffffffffff033bdef4000000c6319ffffffffffffffff"),
                (x"fffffffffffffff0318c6301fffc006318cfffffffffffffff"),
                (x"ffffffffffffffff818c65980fffffffffffffffffffffffff"),

                -- 2_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"ffffffffffffffffd6b5ad6b573ab5ad6ae77fffffffffffff"),
                (x"fffffffffffffeead6a845ef5ad517ba108ab9ceffffffffff"),
                (x"fffffffffffb9d545ef7ba117422f7bdef7422b577ffffffff"),
                (x"fffffffffffb9d545ef7ba117422f7bdef7422b577ffffffff"),
                (x"fffffffffffd6a84210845ee8422f7456b542108afffffffff"),
                (x"ffffffffff756b545ef7ba11742115aa117ba108abbfffffff"),
                (x"ffffffffff756b5ad6a845dd5422a8bdee8456b5abbfffffff"),
                (x"ffffffffff756b5ad6a845dd5422a8bdee8456b5abbfffffff"),
                (x"fffffffffdad6a8455c94dd2ead5c9ba52eaa2b5ad5dffffff"),
                (x"fffffffffdaa108bb937bdef7bdef7bdee972108755dffffff"),
                (x"ffffffffee456b7abaf7bdef7bdef7bdef775508756ae77fff"),
                (x"ffffffffee439d7abaf7bdef7bdef7bdef7756f773aae77fff"),
                (x"fffffff7aeaf7a87258c632f7bdef76318c4baf7ebaae777ff"),
                (x"fffffff7aeaf7a87258c632f7bdef76318c4baf7ebaae777ff"),
                (x"fffffff7b57252875ca0002f7bdef700005bb9084b9d5af7ff"),
                (x"fffffff7b575ef575c80002f7bdef700004bbab5bbbb5af7ff"),
                (x"fffffff7ae70015edc8739ef7bdef739ce4bf6b50740e777ff"),
                (x"fffffffffd7000e05c9291ef7bdef73ca44b81ce0741de83ff"),
                (x"fffffffffd7000e05c9291ef7bdef73ca44b81ce0741de83ff"),
                (x"fffffffffde801d026f7bdef7bdef7bdef7483bd003e007fff"),
                (x"ffffffffff0000003137bdef7bdef7bdee96000007ffffffff"),
                (x"ffffffffffffff42800c62537bdee94b18029694ffffffffff"),
                (x"fffffffffffd285295c42318c6318c614a421294ffffffffff"),
                (x"fffffffffffd285295c42318c6318c614a421294ffffffffff"),
                (x"ffffffffff75285294242109ef7bc42108e090a5a7ffffffff"),
                (x"fffffffff429084700a10843ef7bc10b9c508484a7ffffffff"),
                (x"ffffffffee214a5280a42043ef7bc10908520421253fffffff"),
                (x"fffffffff46108e004052909ef7bc4214a021021253fffffff"),
                (x"fffffffff46108e004052909ef7bc4214a021021253fffffff"),
                (x"ffffffffe04b180f80a42049ef7bc40908021084703fffffff"),
                (x"ffffffffff0001ff80810849ef7bc421080239ce283fffffff"),
                (x"ffffffffffffffff81c42109def7bd239c0026f707ffffffff"),
                (x"fffffffffffffffffc0e757deef7bdef7bff8000ffffffffff"),
                (x"fffffffffffffffffc0e757deef7bdef7bff8000ffffffffff"),
                (x"ffffffffffffffffffe00747eef40c67ffffffffffffffffff"),
                (x"ffffffffffffffffffe0033dd6300007ffffffffffffffffff"),
                (x"ffffffffffffffffffe0032d66301fffffffffffffffffffff"),

                -- 2_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffb9ce756b5ad5ce739dffffffffffffffff"),
                (x"fffffffffffffee75515ad517bdee8456ae77fffffffffffff"),
                (x"fffffffffffd6b742117bdef7bdef7ba108abbffffffffffff"),
                (x"ffffffffff75ee8aa2f7ba2b5ad6a842115455ceffffffffff"),
                (x"ffffffffff75ee8aa2f7ba2b5ad6a842115455ceffffffffff"),
                (x"ffffffffffadef545d15ad51742115aa108aa2b577ffffffff"),
                (x"ffffffffeeab9d5ad5c94a6a8bdd08456a8456b577ffffffff"),
                (x"ffffffffeeaa52e726f7bdd354211542115422b5abbfffffff"),
                (x"ffffffffeeaa52e726f7bdd354211542115422b5abbfffffff"),
                (x"ffffffffeeaa537bdef7bdef5422f5aa108aa108abbfffffff"),
                (x"ffffffffff72537bdef7bdee9ad6e8756a8ad508ad5dffffff"),
                (x"ffffffffffeb197bdef7bdef7ad6e8739d543ab5455dffffff"),
                (x"fffffffffff8017bdd8c63137ad508739d543ab5456bdeffff"),
                (x"fffffffffff8017bdc0001537ad515739cead5ceababdeffff"),
                (x"fffffffffff8017bdc0001537ad515739cead5ceababdeffff"),
                (x"fffffffffff8017bdc000113773915bb9dd755ceababdeffff"),
                (x"fffffffffff8017bdce7392f77390e4f7bded5ce73bbffffff"),
                (x"fffffffffff8017bdcf2912f773aaea77aeed5ceebbbffffff"),
                (x"fffffffffff8017bdef7bdef74a5ceef7aeebbbda77fffffff"),
                (x"fffffffffff8017bdef7bdef74a5ceef7aeebbbda77fffffff"),
                (x"fffffffffff8009bdef7bdef74a5d4ef7aeef694ffffffffff"),
                (x"fffffffffffffe04def7bdee963294a529da7fffffffffffff"),
                (x"fffffffffffffff0018c6318ca50a5a529ffffffffffffffff"),
                (x"ffffffffffffffffd3c529084210242d29ffffffffffffffff"),
                (x"ffffffffffffffffd3c529084210242d29ffffffffffffffff"),
                (x"ffffffffffffffffd3c10848508424294b4fffffffffffffff"),
                (x"fffffffffffffffa7bc5294a408484294b4fffffffffffffff"),
                (x"fffffffffffffffa7bc4210a429485714b4fffffffffffffff"),
                (x"fffffffffffffffa7bc1090a408424a14a5a7fffffffffffff"),
                (x"fffffffffffffffa7bc1090a408424a14a5a7fffffffffffff"),
                (x"fffffffffffffffa7bc1091c108494a14a577fffffffffffff"),
                (x"fffffffffffffffa7bc10869408424a108eeffffffffffffff"),
                (x"fffffffffffffffff7a1092974a68e277bdeffffffffffffff"),
                (x"fffffffffffffffff7bdef6b5739dd6319d07fffffffffffff"),
                (x"fffffffffffffffff7bdef6b5739dd6319d07fffffffffffff"),
                (x"fffffffffffffffffd8c630000001def7ac07fffffffffffff"),
                (x"ffffffffffffffffb18c6001fffc0c6318c07fffffffffffff"),
                (x"fffffffffffffffffffffffff0019663180fffffffffffffff"),

                -- 2_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce739dffffffffffffffff"),
                (x"ffffffffffffffffd6b5ad6b573ab5756b577fffffffffffff"),
                (x"fffffffffffffeead517bd6a8ad515aa108ad5ceffffffffff"),
                (x"fffffffffffb9d5422a845eb74211542115aa2b577ffffffff"),
                (x"fffffffffffb9d5422a845eb74211542115aa2b577ffffffff"),
                (x"fffffffffffd6a8ba115add17422a8456a842108afffffffff"),
                (x"ffffffffff72117ba10842108422a842108422f7abbfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d08abbfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d08abbfffffff"),
                (x"fffffffffdadef7422f7bdd17bdd17bdef7ba2b5ad7bffffff"),
                (x"fffffffffd45ee84210845ef7bdef7bdee842108ad7bffffff"),
                (x"fffffff7ae42108421084211742108ba10842108ad7bffffff"),
                (x"fffffff7b5456a8421084210842108456a842108ad5dffffff"),
                (x"fffffeb9c8456a8421084210842108456a8422b5455ddeffff"),
                (x"fffffeb9c8456a8421084210842108456a8422b5455ddeffff"),
                (x"fffff756a8aa108aa2a84210842108456a8422b5455ddeffff"),
                (x"fffff756a872115422a84210842108ad6a8aa1ce439ddeffff"),
                (x"fffffeb9c8756b5421c84551542108756a8ad5ceab9ddeffff"),
                (x"fffffff7b5ed6ae457a84550e42115756a8abab5abbbffffff"),
                (x"fffffff7b5ed6ae457a84550e42115756a8abab5abbbffffff"),
                (x"ffffffffe0ef7ae43bb5ab90e42115739d5abab573bbffffff"),
                (x"ffffffffffffffde97ae776bdad6aeeb9d5775ce777fffffff"),
                (x"ffffffffffffff4290bdef7a573bbd2f7aee93bdefffffffff"),
                (x"fffffffffffffe5210a529084210842108e29084a7ffffffff"),
                (x"fffffffffffffe5210a529084210842108e29084a7ffffffff"),
                (x"fffffffffffd28421094a38810842109084a14a5253fffffff"),
                (x"fffffffffffb9c4090b4a1485294a529085a3884291dffffff"),
                (x"ffffffffffa5285211d4a14842108421085050a52381ffffff"),
                (x"ffffffffff0108129014a10810842109084a01ce6781ffffff"),
                (x"ffffffffff0108129014a10810842109084a01ce6781ffffff"),
                (x"ffffffffff0318c091c529021084210842470000603fffffff"),
                (x"ffffffffff03189603ae73881213def108477fffffffffffff"),
                (x"fffffffffff800007c1def7bd0018c67bde07fffffffffffff"),
                (x"ffffffffffffffffffe003180003a31f7a0fffffffffffffff"),
                (x"ffffffffffffffffffe003180003a31f7a0fffffffffffffff"),
                (x"ffffffffffffffffffe0031800019eeb19ffffffffffffffff"),
                (x"fffffffffffffffffffff800000196b318cfffffffffffffff"),
                (x"fffffffffffffffffffffffff0018c63180fffffffffffffff"),

                -- 2_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffdce739d5ad6b5739cefffffffffffffff"),
                (x"fffffffffffffff73aa8422f7bdd15aa11573bffffffffffff"),
                (x"fffffffffffffeeaa117bdef7bdef7ba10845eb5ffffffffff"),
                (x"fffffffffffb9d545508422b5ad6a8bdee8aa2f777ffffffff"),
                (x"fffffffffffb9d545508422b5ad6a8bdee8aa2f777ffffffff"),
                (x"ffffffffff756a8aa115ad508bdd15aa117456f7afffffffff"),
                (x"ffffffffff756b5422a842117422a94b9d5ad5ceabbfffffff"),
                (x"ffffffffff756b54210845508ad537bdee973929abbfffffff"),
                (x"ffffffffff756b54210845508ad537bdee973929abbfffffff"),
                (x"ffffffffeead6b545508456e8ad6f7bdef7bdd29abbfffffff"),
                (x"ffffffffeead6a845515aa2f54a6f7bdef7bdd2977ffffffff"),
                (x"ffffffffeeab9c845515aa2f5bdef7bdef7bdd8cefffffffff"),
                (x"ffffffffeeab9c8ab90e72115bdd2c63197bdc00ffffffffff"),
                (x"fffffffffdab9c8abaae75515bdd2500017bdc00ffffffffff"),
                (x"fffffffffdab9c8abaae75515bdd2500017bdc00ffffffffff"),
                (x"fffffffffdab9c8ab9d7bd50ebdd2400017bdc00ffffffffff"),
                (x"fffffffffd777b5ab9c94b90ebdee439cf7bdc00ffffffffff"),
                (x"fffffffffd777b5ab9d4a3aaebdee491cf7bdc00ffffffffff"),
                (x"ffffffffffef7aeaf5ddeb9c9bdef7bdef7bdc00ffffffffff"),
                (x"ffffffffffef7aeaf5ddeb9c9bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffffd29d775dded1c9bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffa7694a528c4a6f7bdef7483ffffffffffff"),
                (x"ffffffffffffffffd0a52d1c56318c6318007fffffffffffff"),
                (x"fffffffffffffffa14810948521294a528e253ffffffffffff"),
                (x"fffffffffffffffa14810948521294a528e253ffffffffffff"),
                (x"fffffffffffffffa1081090a4084a4a7bc12d3ffffffffffff"),
                (x"fffffffffffffff71484210a40842ea7bd429694ffffffffff"),
                (x"ffffffffffffff42902e750810848ea7bd42ba94ffffffffff"),
                (x"ffffffffffffff4714a528084210a4a7bdea1484ffffffffff"),
                (x"ffffffffffffff4714a528084210a4a7bdea1484ffffffffff"),
                (x"ffffffffffffff4a102e70081084a1a7bdea1000ffffffffff"),
                (x"fffffffffffffe0631800388408425efbdea5c00ffffffffff"),
                (x"fffffffffffffff026e0076b5ef7def77a0003ffffffffffff"),
                (x"fffffffffffffff0001def7bdef7bdef7a0fffffffffffffff"),
                (x"fffffffffffffff0001def7bdef7bdef7a0fffffffffffffff"),
                (x"fffffffffffffff0318000000ef7c36001ffffffffffffffff"),
                (x"fffffffffffffff0318c603e0633be63180fffffffffffffff"),
                (x"fffffffffffffffffffffffff00196b3180fffffffffffffff"),

                -- 2_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"ffffffffffffffffd6b5ad6b573ab5ad6ae77fffffffffffff"),
                (x"fffffffffffffeead6a845ef5ad517ba108ab9ceffffffffff"),
                (x"fffffffffffb9d545ef7ba117422f7bdef7422b577ffffffff"),
                (x"fffffffffffb9d545ef7ba117422f7bdef7422b577ffffffff"),
                (x"fffffffffffd6a84210845ee8422f7456b542108afffffffff"),
                (x"ffffffffff756b545ef7ba11742115aa117ba108abbfffffff"),
                (x"ffffffffff756b5ad6a845dd5422a8bdee8456b5abbfffffff"),
                (x"ffffffffff756b5ad6a845dd5422a8bdee8456b5abbfffffff"),
                (x"fffffffffdad6a8455c94dd2ead5c9ba52eaa2b5abbbffffff"),
                (x"fffffffffdaa108bb937bdef7bdef7bdee972108ad7bffffff"),
                (x"ffffffb9d5ab9c8abaf7bdef7bdef7bdef7756f7ad5dffffff"),
                (x"ffffffb9d5739d7abaf7bdef7bdef7bdef7756f7755ddeffff"),
                (x"fffffeb9d5777b77258c632f7bdef76318c4b908ed5ddeffff"),
                (x"fffffeb9d5777b77258c632f7bdef76318c4b908ed5ddeffff"),
                (x"fffffed6ae7252875ca0002f7bdef700005bb9084b9ddeffff"),
                (x"fffffed6bd75ef575c80002f7bdef700004bbab5bf5ddeffff"),
                (x"fffffeb9dde8015edc8739ef7bdef739ce4bf6b503bbffffff"),
                (x"fffff077a0e800e05c9291ef7bdef73ca44b81ce03bbffffff"),
                (x"fffff077a0e800e05c9291ef7bdef73ca44b81ce03bbffffff"),
                (x"ffffff801fe801d026f7bdef7bdef7bdef7483bd077fffffff"),
                (x"ffffffffff07fe003137bdef7bdef7bdee96000007ffffffff"),
                (x"ffffffffffffff42940c62537bdee94b18001694ffffffffff"),
                (x"ffffffffffffff4210852b18c6318c6108e294a5a7ffffffff"),
                (x"ffffffffffffff4210852b18c6318c6108e294a5a7ffffffff"),
                (x"fffffffffffd285205c10909ef7bc421081294a5a3bfffffff"),
                (x"fffffffffffd284084ae7043ef7bc108425038842169ffffff"),
                (x"ffffffffffa1081090a42043ef7bc109085014a5291dffffff"),
                (x"ffffffffffa1081210052909ef7bc4214a0081ce2329ffffff"),
                (x"ffffffffffa1081210052909ef7bc4214a0081ce2329ffffff"),
                (x"ffffffffff039c4210042049ef7bc40908507c006241ffffff"),
                (x"ffffffffff014ae710042109ef7bc40842407fff003fffffff"),
                (x"fffffffffff80174800e713bdef7a42108e07fffffffffffff"),
                (x"fffffffffffffe007ffdef7bdf7bdeab9c0fffffffffffffff"),
                (x"fffffffffffffe007ffdef7bdf7bdeab9c0fffffffffffffff"),
                (x"fffffffffffffffffffffb180ef7c3e801ffffffffffffffff"),
                (x"fffffffffffffffffffff8000633be6001ffffffffffffffff"),
                (x"fffffffffffffffffffffffe0632d66001ffffffffffffffff"),

                -- 2_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffb9ce756b5ad5ce739dffffffffffffffff"),
                (x"fffffffffffffee75515ad517bdee8456ae77fffffffffffff"),
                (x"fffffffffffd6b742117bdef7bdef7ba108abbffffffffffff"),
                (x"ffffffffff75ee8aa2f7ba2b5ad6a842115455ceffffffffff"),
                (x"ffffffffff75ee8aa2f7ba2b5ad6a842115455ceffffffffff"),
                (x"ffffffffffadef545d15ad51742115aa108aa2b577ffffffff"),
                (x"ffffffffeeab9d5ad5c94a6a8bdd08456a8456b577ffffffff"),
                (x"ffffffffeeaa52e726f7bdd354211542108456b577ffffffff"),
                (x"ffffffffeeaa52e726f7bdd354211542108456b577ffffffff"),
                (x"ffffffffeeaa537bdef7bdef5422f542115456b5abbfffffff"),
                (x"ffffffffff72537bdef7bdee9ad6e8aa115422b5abbfffffff"),
                (x"ffffffffffeb197bdef7bdef7ad6e8aa115421ceabbfffffff"),
                (x"fffffffffff8017bdd8c63137ad5087210eaa1ceabbfffffff"),
                (x"fffffffffff8017bdc0001537ad515756aeaa1ceaf7fffffff"),
                (x"fffffffffff8017bdc0001537ad515756aeaa1ceaf7fffffff"),
                (x"fffffffffff8017bdc000113773915bb9ceaa1ceaf7fffffff"),
                (x"fffffffffff8017bdce7392f77390e4b9cead7bd777fffffff"),
                (x"fffffffffff8017bdcf2912f773aaea39cead7bd777fffffff"),
                (x"fffffffffff8017bdef7bdef74a5ceeb9ddabbbdefffffffff"),
                (x"fffffffffff8017bdef7bdef74a5ceeb9ddabbbdefffffffff"),
                (x"fffffffffff8009bdef7bdef74a5d4eb9dd77694ffffffffff"),
                (x"fffffffffffffe04def7bdee963294a529da7fffffffffffff"),
                (x"fffffffffffffff0018c6318c295d4294b4fffffffffffffff"),
                (x"ffffffffffffff423a94a52842948509085a7fffffffffffff"),
                (x"ffffffffffffff423a94a52842948509085a7fffffffffffff"),
                (x"ffffffffffffff4287d4a10a1210a409084a7fffffffffffff"),
                (x"fffffffffffd2852d3d4a3821210a42108577fffffffffffff"),
                (x"fffffffffffd28e2d3d4a388108494704242d3ffffffffffff"),
                (x"fffffffffff9085a7bd4a10a421080294a5753ffffffffffff"),
                (x"fffffffffff9085a7bd4a10a421080294a5753ffffffffffff"),
                (x"fffffffffff8004a7bd4a04a10848070424a53ffffffffffff"),
                (x"fffffffffff8017a7bdde94212108e0318c603ffffffffffff"),
                (x"fffffffffffffe0003bef7bdd2109d05ee907fffffffffffff"),
                (x"ffffffffffffffff83bdef7bdef7bde800007fffffffffffff"),
                (x"ffffffffffffffff83bdef7bdef7bde800007fffffffffffff"),
                (x"fffffffffffffffffc0c60fdd000000318c07fffffffffffff"),
                (x"ffffffffffffffff818c67bac003e06318c07fffffffffffff"),
                (x"ffffffffffffffff8196b5980fffffffffffffffffffffffff"),

                -- 3_character_0_0
                (x"fffffffffffffffffffef7bdef7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffffffef7bdef7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffffbc739ce739ce739cfef7fffffffffffff"),
                (x"ffffffffffffffff1ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffff438c6318c6318c6318c6739e94ffffffffff"),
                (x"fffffffffffd29e18c6318c6318c6318c6339fdea7ffffffff"),
                (x"fffffffffffd29e18c6318c6318c6318c6339fdea7ffffffff"),
                (x"fffffffffffd28718c6318c6318c6318c6339ce7a7ffffffff"),
                (x"ffffffffffa7bc318ce318c6318c6318c6739ce7f53fffffff"),
                (x"ffffffffffa1ce318ce738c6318c6319ce739ce7f53fffffff"),
                (x"ffffffffffa1ce318ce738c6318c6319ce739ce7f53fffffff"),
                (x"ffffffffffa0c6718ce739ce739ce739ce739ce7f53fffffff"),
                (x"ffffffffffa0c7e18ce739ce739ce739ce739fdef53fffffff"),
                (x"ffffffffffa1cfe18ce739ce739ce739ce739fdef53fffffff"),
                (x"ffffffffffa7bde38c7ef1ce739ce73fbc739fdef53fffffff"),
                (x"ffffffffffa7bdef1c7ef1ce739ce7f7bc73fbdef53fffffff"),
                (x"ffffffffffa7bdef1c7ef1ce739ce7f7bc73fbdef53fffffff"),
                (x"fffffffffffd29ef1ce73f8e739ce7f1ce73fbdea53fffffff"),
                (x"fffffffffffd29ef78e73fbc739cfef1ce7f7bdea7ffffffff"),
                (x"ffffffffffffff4f7bc739e9ef7bd439cfef7a94ffffffffff"),
                (x"fffffffffffffffa7bdef7a94a53d4f7bdef53ffffffffffff"),
                (x"fffffffffffffffa7bdef7a94a53d4f7bdef53ffffffffffff"),
                (x"ffffffffffffff43d29ef1fc718cfe3fbd4a1e94ffffffffff"),
                (x"fffffffffffd2871fa9defbb4a529405294f0ce7a7ffffffff"),
                (x"ffffffffffa7bc33fa9defbdef7bdef77bdf1c63f53fffffff"),
                (x"fffffffff4a7bc7f7a9defbdef7bdef7bd4f78e7f529ffffff"),
                (x"fffffffff4a7bc7f7a9defbdef7bdef7bd4f78e7f529ffffff"),
                (x"fffffffff4f5294a7a94a77d4f7a9ef77b4f5294a7a9ffffff"),
                (x"fffffffffda7bdea0294a529def7b4a5294053def53bffffff"),
                (x"fffffffff4ed28000294a77bdef7bded29400000a769ffffff"),
                (x"fffffffff4a5294a029ef1c67f78e33fbd405294a529ffffff"),
                (x"fffffffff4a5294a029ef1c67f78e33fbd405294a529ffffff"),
                (x"ffffffffffa529400294a78fea53c7f529400294a53fffffff"),
                (x"ffffffffffffffffd3c73d28000014a1cfea7fffffffffffff"),
                (x"ffffffffffffffffd29ef0cfea53c71fbd4a7fffffffffffff"),
                (x"ffffffffffffffff8294a529400294a529407fffffffffffff"),
                (x"ffffffffffffffff8294a529400294a529407fffffffffffff"),
                (x"fffffffffffffffffc1ef7a9400294f7bc0fffffffffffffff"),
                (x"fffffffffffffffffc14a7a80ffc14f5280fffffffffffffff"),
                (x"fffffffffffffffffc1ef1fc0ffc1e3fbc0fffffffffffffff"),

                -- 3_character_0_1
                (x"fffffffffffffffffe94a5294f7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffffe94a5294f7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffa53def1c6318c6339cfef7fffffffffffff"),
                (x"ffffffffffffff4f1ce739ce739c6318c633fbffffffffffff"),
                (x"fffffffffffd29e39ce739ce318c631fbcf1bfdeffffffffff"),
                (x"fffffffffffd28739ce738c6318c63f0c63295efffffffffff"),
                (x"fffffffffffd28739ce738c6318c63f0c63295efffffffffff"),
                (x"ffffffffffa7bc73f8e318cfef78fe1bdfe1d0a5a7ffffffff"),
                (x"ffffffffffa7bc7f78e73fbc7f7bc37fbc0180a5a7ffffffff"),
                (x"fffffffff4f7bdef1cfef7a9418c7ef528078063a7ffffffff"),
                (x"fffffffff4f7bdef1cfef7a9418c7ef528078063a7ffffffff"),
                (x"fffffffff4f7bdef1fd4a51e37bfdef5280781efa7ffffffff"),
                (x"fffffffff4f7bdef780f7bfdef7bdef7bd4f51ef07ffffffff"),
                (x"fffffffff4f7bdef501ef7bdef7a800001ef7800ffffffffff"),
                (x"ffffffffffa7bdef7814a7bdea50190000000000ffffffffff"),
                (x"ffffffffffa7bdea7bd4a0294a5019ce72739c00ffffffffff"),
                (x"ffffffffffa7bdea7bd4a0294a5019ce72739c00ffffffffff"),
                (x"fffffffffffd29ea7a94a02947bc199ce6739c00ffffffffff"),
                (x"fffffffffffd294a5294a0294f79fe9d28329463ffffffffff"),
                (x"ffffffffffffffea5294a0294f7bcfa0c6f780a5a7ffffffff"),
                (x"fffffffffffffffa5294a0294f7bdea3de078063a7ffffffff"),
                (x"fffffffffffffffa5294a0294f7bdea3de078063a7ffffffff"),
                (x"fffffffffffffffffe94a5014a53dea3df478000ffffffffff"),
                (x"fffffffffffffffffc14a528000014a5294003ffffffffffff"),
                (x"ffffffffffffffff83c73d29da5294a5280fffffffffffffff"),
                (x"ffffffffffffffffd0631fa9df7bbe3fbd4fffffffffffffff"),
                (x"ffffffffffffffffd0631fa9df7bbe3fbd4fffffffffffffff"),
                (x"fffffffffffffff078fef1c67a528739cfefffffffffffffff"),
                (x"fffffffffffffff07a8738fb400014f7bd4fffffffffffffff"),
                (x"fffffffffffffff052873f69e18fc0a5280fffffffffffffff"),
                (x"ffffffffffffffff829ef768739fc0ed280fffffffffffffff"),
                (x"ffffffffffffffff829ef768739fc0ed280fffffffffffffff"),
                (x"ffffffffffffffff8014a529ef7a8019cf4fffffffffffffff"),
                (x"ffffffffffffffff8280052940001e3d294fffffffffffffff"),
                (x"fffffffffffffffffc14a0000a5294f529ffffffffffffffff"),
                (x"ffffffffffffffffffe0053c718cfea7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0053c718cfea7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0053def7a9407ffffffffffffffffff"),
                (x"fffffffffffffffffffffd294a5280ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83de39fc0ffffffffffffffffffff"),

                -- 3_character_0_2
                (x"ffffffffffffffffffffffbdea5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffffffbdea5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffdef78e739ce7f7bd4a7fffffffffffff"),
                (x"fffffffffffffffa78e738c6318c6318c67f53ffffffffffff"),
                (x"ffffffffffffff4f1c6318c6318c6318c633fa94ffffffffff"),
                (x"fffffffffffd29e38c6319cfef7bc739ce319fdea7ffffffff"),
                (x"fffffffffffd29e38c6319cfef7bc739ce319fdea7ffffffff"),
                (x"fffffffffffd28719ce73f9e5294aff7bde39fdea7ffffffff"),
                (x"ffffffffffa7bc339cef794a3a53c51bdfef7bdef53fffffff"),
                (x"ffffffffffa7bc3f1de52be83003d478c6ff7a94f53fffffff"),
                (x"ffffffffffa7bc3f1de52be83003d478c6ff7a94f53fffffff"),
                (x"ffffffffffa1cfe3bcaf78c03003c07fbc37fa94f53fffffff"),
                (x"ffffffffffa1cf4f15e318c03a53c07fbde1fa94a53fffffff"),
                (x"ffffffffffa000f7d3cf78e83a53d47fbdea3def053fffffff"),
                (x"ffffffffffa001ef001ef3c637bfcff7bc007bde053fffffff"),
                (x"ffffffffffa5294f032000294a52940001907a94a53fffffff"),
                (x"ffffffffffa5294f032000294a52940001907a94a53fffffff"),
                (x"ffffffffffa5280a0339ce4e739ce7ce73905000a53fffffff"),
                (x"fffffffffff8000a53339cfd4a529e9ce79a500007ffffffff"),
                (x"fffffffffffffe0f53339f8a5294a3f4e79a7800ffffffffff"),
                (x"fffffffffffffe0a7874a1463003cf1d28ff5000ffffffffff"),
                (x"fffffffffffffe0a7874a1463003cf1d28ff5000ffffffffff"),
                (x"fffffffffffd29ea79f4a3c03003c0f528ff53dea7ffffffff"),
                (x"fffffffff4a7bc33d3d4a3e83003d4f529ea1c63f529ffffff"),
                (x"ffffffd28719ce7f5294a51eff7bdea5294a78e738cf4a7fff"),
                (x"fffffa1cfea5294a529defa94a5294f77b4a5294a53c73d3ff"),
                (x"fffffa1cfea5294a529defa94a5294f77b4a5294a53c73d3ff"),
                (x"fffffa1cf4ef7b4a53dde9ce739ce73f7bea5294ef6873d3ff"),
                (x"fffff0529da5294a0294a7bdef7bdef529405294a53b4a03ff"),
                (x"ffffff8014a0c67a0294a5294a5294a5294050e71d28007fff"),
                (x"ffffffffe0f1ce7a0294a53bdef7bda5294050e73f80007fff"),
                (x"ffffffffe0f1ce7a0294a53bdef7bda5294050e73f80007fff"),
                (x"ffffffffe0a7bde00294a78e318c67f5294003def501ffffff"),
                (x"ffffffffff00000f8014a53c739cfea528007c00003fffffff"),
                (x"ffffffffffffffffd3c73d29400294a1cfea7fffffffffffff"),
                (x"ffffffffffffffff829ef0cf4002871fbd407fffffffffffff"),
                (x"ffffffffffffffff829ef0cf4002871fbd407fffffffffffff"),
                (x"ffffffffffffffff8294a528000014a529407fffffffffffff"),
                (x"fffffffffffffffffc1ef0fc0ffc1e1fbc0fffffffffffffff"),
                (x"fffffffffffffffffc14a5280ffc14a5280fffffffffffffff"),

                -- 3_character_0_3
                (x"ffffffffffffffffffdef7bdea5294a529ffffffffffffffff"),
                (x"ffffffffffffffffffdef7bdea5294a529ffffffffffffffff"),
                (x"ffffffffffffffff78e738c6318c67f7bd4a7fffffffffffff"),
                (x"ffffffffffffffe38c6318c6739ce739ce7f53ffffffffffff"),
                (x"ffffffffffffbcf1bfc318c6318ce739ce73fa94ffffffffff"),
                (x"fffffffffffbde528c7ef0c6318c6339ce739e94ffffffffff"),
                (x"fffffffffffbde528c7ef0c6318c6339ce739e94ffffffffff"),
                (x"ffffffffffa14b41f9e31f8fef78e319cfe39fdea7ffffffff"),
                (x"ffffffffffa14a0183cf78fde39fde39cfef1fdea7ffffffff"),
                (x"ffffffffffa0c607829ef7863a529ef1ce7f7bdef53fffffff"),
                (x"ffffffffffa0c607829ef7863a529ef1ce7f7bdef53fffffff"),
                (x"ffffffffffa3de07829ef7bcf18df4a7bc7f7bdef53fffffff"),
                (x"ffffffffff03df4f53def7bdef7bcf7801ef7bdef53fffffff"),
                (x"fffffffffff801ef78000029ef7bdef0014f7bdef53fffffff"),
                (x"fffffffffff80000000006414f7bdea001ef7bdea7ffffffff"),
                (x"fffffffffff800739f39ce414a5280a7bdea7bdea7ffffffff"),
                (x"fffffffffff800739f39ce414a5280a7bdea7bdea7ffffffff"),
                (x"fffffffffff800739e739e40fa5280a529ea7a94ffffffffff"),
                (x"fffffffffff8c6528e939f9fea5280a5294a5294ffffffffff"),
                (x"ffffffffffa14a07bc74a3fdea5280a5294a7bffffffffffff"),
                (x"ffffffffffa0c60781f4a7bdea5280a5294fffffffffffffff"),
                (x"ffffffffffa0c60781f4a7bdea5280a5294fffffffffffffff"),
                (x"fffffffffff80007d1f4a7bd4a5014a529ffffffffffffffff"),
                (x"fffffffffffffe005294a500000294a001ffffffffffffffff"),
                (x"ffffffffffffffff8294a5294ef6943fbc0fffffffffffffff"),
                (x"ffffffffffffffffd3c73fbbeef69e18c74fffffffffffffff"),
                (x"ffffffffffffffffd3c73fbbeef69e18c74fffffffffffffff"),
                (x"fffffffffffffffff8e739e9439c67f1cfe07fffffffffffff"),
                (x"ffffffffffffffffd3def5000a53a33d29e07fffffffffffff"),
                (x"ffffffffffffffff8294a03c3f7a9d3d29407fffffffffffff"),
                (x"ffffffffffffffff829de83c739e9df5280fffffffffffffff"),
                (x"ffffffffffffffff829de83c739e9df5280fffffffffffffff"),
                (x"ffffffffffffffffd0e31829ef7a94a0000fffffffffffffff"),
                (x"ffffffffffffffffd2873f800a529405280fffffffffffffff"),
                (x"fffffffffffffffffe9ef529400000a001ffffffffffffffff"),
                (x"fffffffffffffffffff4a78e339fd407ffffffffffffffffff"),
                (x"fffffffffffffffffff4a78e339fd407ffffffffffffffffff"),
                (x"ffffffffffffffffffe00529ef7bd407ffffffffffffffffff"),
                (x"fffffffffffffffffffff8294a5294ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83c7f7bc0ffffffffffffffffffff"),

                -- 3_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffef7bdef7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffffbc739ce739ce739cfef7fffffffffffff"),
                (x"ffffffffffffffff1ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffff438c6318c6318c6318c6739e94ffffffffff"),
                (x"ffffffffffffff438c6318c6318c6318c6739e94ffffffffff"),
                (x"fffffffffffd29e18c6318c6318c6318c6339fdea7ffffffff"),
                (x"fffffffffffd28718c6318c6318c6318c6339ce7a7ffffffff"),
                (x"ffffffffffa7bc318ce318c6318c6318c6739ce7f53fffffff"),
                (x"ffffffffffa7bc318ce318c6318c6318c6739ce7f53fffffff"),
                (x"ffffffffffa1ce318ce738c6318c6319ce739ce7f53fffffff"),
                (x"ffffffffffa0c6718ce739ce739ce739ce739ce7f53fffffff"),
                (x"ffffffffffa0c7e18ce739ce739ce739ce739fdef53fffffff"),
                (x"ffffffffffa1cfe18ce739ce739ce739ce739fdef53fffffff"),
                (x"ffffffffffa7bde38c7ef1ce739ce73fbc739fdef53fffffff"),
                (x"ffffffffffa7bde38c7ef1ce739ce73fbc739fdef53fffffff"),
                (x"ffffffffffa7bdef1c7ef1ce739ce7f7bc73fbdef53fffffff"),
                (x"fffffffffffd29ef1ce73f8e739ce7f1ce73fbdea53fffffff"),
                (x"fffffffffffd29ef78e73fbc739cfef1ce7f7bdea7ffffffff"),
                (x"ffffffffffffff4f7bc739e9ef7bd439cfef7a94ffffffffff"),
                (x"ffffffffffffff4f7bc739e9ef7bd439cfef7a94ffffffffff"),
                (x"fffffffffffffffa7bdef7a94a53d4f7bdef53ffffffffffff"),
                (x"ffffffffffffff4f529defbb4a529405294a53ffffffffffff"),
                (x"fffffffffffd29e3fa9defbde18fdef77bdf7a94ffffffffff"),
                (x"ffffffffffa7bc7f7a9defbdef7bdef7bd4f1e94ffffffffff"),
                (x"ffffffffffa7bc7f7a9defbdef7bdef7bd4f1e94ffffffffff"),
                (x"fffffffff4a529ea7a94a77d4f7bdef77b4f7a94a7ffffffff"),
                (x"fffffffff4a7bdea7a94a529def7b4a5294f5294a53fffffff"),
                (x"ffffffffffa5294003d4a5294a5294a001ea53dea53fffffff"),
                (x"ffffffffffa529da5294a77bdef694a001ef7bbda03fffffff"),
                (x"ffffffffffa529da5294a77bdef694a001ef7bbda03fffffff"),
                (x"fffffffffffd294a03c738cfea53c7f5294ef694a7ffffffff"),
                (x"fffffffffffffe00029ef7a800029ea5280a529407ffffffff"),
                (x"fffffffffffffffffc14a1cfe00294a5280003ffffffffffff"),
                (x"fffffffffffffffffc1ef7a94f7814a001ffffffffffffffff"),
                (x"fffffffffffffffffc1ef7a94f7814a001ffffffffffffffff"),
                (x"ffffffffffffffffffe0050e7f780007ffffffffffffffffff"),
                (x"fffffffffffffffffffff83d4a501fffffffffffffffffffff"),
                (x"fffffffffffffffffffff8294a501fffffffffffffffffffff"),

                -- 3_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294f7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffa53def1c6318c6339cfef7fffffffffffff"),
                (x"ffffffffffffff4f1ce739ce739c6318c633fbffffffffffff"),
                (x"fffffffffffd29e39ce739ce318c631fbcf1bfdeffffffffff"),
                (x"fffffffffffd29e39ce739ce318c631fbcf1bfdeffffffffff"),
                (x"fffffffffffd28739ce738c6318c63f0c63295efffffffffff"),
                (x"ffffffffffa7bc73f8e318cfef78fe1bdfe1d0a5a7ffffffff"),
                (x"ffffffffffa7bc7f78e73fbc7f7bc37fbc0180a5a7ffffffff"),
                (x"ffffffffffa7bc7f78e73fbc7f7bc37fbc0180a5a7ffffffff"),
                (x"fffffffff4f7bdef1cfef7a9418c7ef528078063a7ffffffff"),
                (x"fffffffff4f7bdef1fd4a51e37bfdef5280781efa7ffffffff"),
                (x"fffffffff4f7bdef780f7bfdef7bdef7bd4f51ef07ffffffff"),
                (x"fffffffff4f7bdef501ef7bdef7a800001ef7800ffffffffff"),
                (x"ffffffffffa7bdef7814a7bdea50190000000000ffffffffff"),
                (x"ffffffffffa7bdef7814a7bdea50190000000000ffffffffff"),
                (x"ffffffffffa7bdea7bd4a0294a5019ce72739c00ffffffffff"),
                (x"fffffffffffd29ea7a94a02947bc199ce6739c00ffffffffff"),
                (x"fffffffffffd294a5294a0294f79fe9d28329463ffffffffff"),
                (x"ffffffffffffffea5294a0294f7bcfa0c6f780a5a7ffffffff"),
                (x"ffffffffffffffea5294a0294f7bcfa0c6f780a5a7ffffffff"),
                (x"ffffffffffffffffd294a0294f7bdea3de078063a7ffffffff"),
                (x"fffffffffffffffffe94a5014a53dea3df478000ffffffffff"),
                (x"fffffffffffffffffc14a53a000014a5294003ffffffffffff"),
                (x"fffffffffffffffffc1ef1e9df7a94a5294fffffffffffffff"),
                (x"fffffffffffffffffc1ef1e9df7a94a5294fffffffffffffff"),
                (x"ffffffffffffffff83c318fd4a53be3fbd4fffffffffffffff"),
                (x"ffffffffffffffff83c73fa87a529439cf4fffffffffffffff"),
                (x"ffffffffffffffff829ef50feef4fea7bd4fffffffffffffff"),
                (x"fffffffffffffff05014a53d4ef4633fbd4fffffffffffffff"),
                (x"fffffffffffffff05014a53d4ef4633fbd4fffffffffffffff"),
                (x"fffffffffffffff07a80053dda50e3f529ffffffffffffffff"),
                (x"fffffffffffffffa7a94a0294a50000529ffffffffffffffff"),
                (x"fffffffffffffff053c73d00000014a529ffffffffffffffff"),
                (x"fffffffffffffff0529ef1cf40029e3fbdffffffffffffffff"),
                (x"fffffffffffffff0529ef1cf40029e3fbdffffffffffffffff"),
                (x"ffffffffffffffffd294a5280a5294f529ffffffffffffffff"),
                (x"fffffffffffffffffbd4a001fffe9e3fbd4fffffffffffffff"),
                (x"ffffffffffffffffd2873fa80fffffffffffffffffffffffff"),

                -- 3_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffbdea5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffdef78e739ce7f7bd4a7fffffffffffff"),
                (x"fffffffffffffffa78e738c6318c6318c67f53ffffffffffff"),
                (x"ffffffffffffff4f1c6318c6318c6318c633fa94ffffffffff"),
                (x"ffffffffffffff4f1c6318c6318c6318c633fa94ffffffffff"),
                (x"fffffffffffd29e38c6319cfef7bc739ce319fdea7ffffffff"),
                (x"fffffffffffd28719ce73f9e5294aff7bde39fdea7ffffffff"),
                (x"ffffffffffa7bc339cef794a3a53c51bdfef7bdef53fffffff"),
                (x"ffffffffffa7bc339cef794a3a53c51bdfef7bdef53fffffff"),
                (x"ffffffffffa7bc3f1de52be83003d478c6ff7a94f53fffffff"),
                (x"ffffffffffa1cfe3bcaf78c03003c07fbc37fa94f53fffffff"),
                (x"ffffffffffa1cf4f15e318c03a53c07fbde1fa94a53fffffff"),
                (x"ffffffffffa000f7d3cf78e83a53d47fbdea3def053fffffff"),
                (x"ffffffffffa001ef001ef3c637bfcff7bc007bde053fffffff"),
                (x"ffffffffffa001ef001ef3c637bfcff7bc007bde053fffffff"),
                (x"ffffffffffa5294f032000294a52940001907a94a53fffffff"),
                (x"ffffffffffa5280a0339ce4e739ce7ce73905000a53fffffff"),
                (x"fffffffffff8000a53339cfd4a529e9ce79a500007ffffffff"),
                (x"fffffffffffffe0f53339f8a5294a3f4e79a7800ffffffffff"),
                (x"fffffffffffffe0f53339f8a5294a3f4e79a7800ffffffffff"),
                (x"fffffffffffffe0a7874a1463003cf1d28ff5000ffffffffff"),
                (x"fffffffffffd29ea79f4a3c03003c0f528ff53dea7ffffffff"),
                (x"fffffffff4f7bdef53d4a3e83003d4f529ea78e73d3fffffff"),
                (x"ffffffd2873d29ea77d4a51eff7bdea5294ef8e73fa9ffffff"),
                (x"ffffffd2873d29ea77d4a51eff7bdea5294ef8e73fa9ffffff"),
                (x"fffffffbc319cfea53ddefa94a5294efbd4a50e718fdffffff"),
                (x"ffffffd29da529ea03d4a1ce739ce7a7bd4053bdf1c74a7fff"),
                (x"ffffffd294a5294a5294a7bdef7bdef5280a7a94ef8f4a7fff"),
                (x"ffffffd29ef5280f8294a5294a5294a529419fdea53d4a7fff"),
                (x"ffffffd29ef5280f8294a5294a5294a529419fdea53d4a7fff"),
                (x"ffffffd2873fbc0f829ef529def7b4a529439fdea529ffffff"),
                (x"ffffff8007f529ffd294a7bc718c67f5280a7a9407ffffffff"),
                (x"ffffffffe00001ff83c738e94f78fea529400000ffffffffff"),
                (x"fffffffffffffffffe9ef78e3a5014a529ffffffffffffffff"),
                (x"fffffffffffffffffe9ef78e3a5014a529ffffffffffffffff"),
                (x"fffffffffffffffffff4a7bdea5014f001ffffffffffffffff"),
                (x"ffffffffffffffffffe0053d40000007ffffffffffffffffff"),
                (x"fffffffffffffffffffff8067003ffffffffffffffffffffff"),

                -- 3_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffdef7bdea5294a529ffffffffffffffff"),
                (x"ffffffffffffffff78e738c6318c67f7bd4a7fffffffffffff"),
                (x"ffffffffffffffe38c6318c6739ce739ce7f53ffffffffffff"),
                (x"ffffffffffffbcf1bfc318c6318ce739ce73fa94ffffffffff"),
                (x"ffffffffffffbcf1bfc318c6318ce739ce73fa94ffffffffff"),
                (x"fffffffffffbde528c7ef0c6318c6339ce739e94ffffffffff"),
                (x"ffffffffffa14b41f9e31f8fef78e319cfe39fdea7ffffffff"),
                (x"ffffffffffa14a0183cf78fde39fde39cfef1fdea7ffffffff"),
                (x"ffffffffffa14a0183cf78fde39fde39cfef1fdea7ffffffff"),
                (x"ffffffffffa0c607829ef7863a529ef1ce7f7bdef53fffffff"),
                (x"ffffffffffa3de07829ef7bcf18df4a7bc7f7bdef53fffffff"),
                (x"ffffffffff03df4f53def7bdef7bcf7801ef7bdef53fffffff"),
                (x"fffffffffff801ef78000029ef7bdef0014f7bdef53fffffff"),
                (x"fffffffffff80000000006414f7bdea001ef7bdea7ffffffff"),
                (x"fffffffffff80000000006414f7bdea001ef7bdea7ffffffff"),
                (x"fffffffffff800739f39ce414a5280a7bdea7bdea7ffffffff"),
                (x"fffffffffff800739e739e40fa5280a529ea7a94ffffffffff"),
                (x"fffffffffff8c6528e939f9fea5280a5294a5294ffffffffff"),
                (x"ffffffffffa14a07bc74a3fdea5280a5294a7bffffffffffff"),
                (x"ffffffffffa14a07bc74a3fdea5280a5294a7bffffffffffff"),
                (x"ffffffffffa0c60781f4a7bdea5280a5294a7fffffffffffff"),
                (x"fffffffffff80007d1f4a7bd4a5014a529ffffffffffffffff"),
                (x"fffffffffffffe005294a5000003b4a001ffffffffffffffff"),
                (x"ffffffffffffffffd294a529eef687f001ffffffffffffffff"),
                (x"ffffffffffffffffd294a529eef687f001ffffffffffffffff"),
                (x"ffffffffffffffffd3c73fbb4a53c31fbc0fffffffffffffff"),
                (x"ffffffffffffffffd0e73d29439e9e3fbc0fffffffffffffff"),
                (x"ffffffffffffffffd3d4a78fdf78f4f5280fffffffffffffff"),
                (x"ffffffffffffffffd3c738c7da53d4a001407fffffffffffff"),
                (x"ffffffffffffffffd3c738c7da53d4a001407fffffffffffff"),
                (x"fffffffffffffffffe9ef0cf4ef7d40529e07fffffffffffff"),
                (x"fffffffffffffffffe8000014a5280a529ea7fffffffffffff"),
                (x"fffffffffffffffffe94a5000000143fbd407fffffffffffff"),
                (x"ffffffffffffffffffc73fa80a50e7f529407fffffffffffff"),
                (x"ffffffffffffffffffc73fa80a50e7f529407fffffffffffff"),
                (x"fffffffffffffffffe9ef529400294a5294fffffffffffffff"),
                (x"ffffffffffffffffd3c73fa9fffc00a7bdefffffffffffffff"),
                (x"fffffffffffffffffffffffff0029e3d294fffffffffffffff"),

                -- 3_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffef7bdef7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffffbc739ce739ce739cfef7fffffffffffff"),
                (x"ffffffffffffffff1ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffff438c6318c6318c6318c6739e94ffffffffff"),
                (x"ffffffffffffff438c6318c6318c6318c6739e94ffffffffff"),
                (x"fffffffffffd29e18c6318c6318c6318c6339fdea7ffffffff"),
                (x"fffffffffffd28718c6318c6318c6318c6339ce7a7ffffffff"),
                (x"ffffffffffa7bc318ce318c6318c6318c6739ce7f53fffffff"),
                (x"ffffffffffa7bc318ce318c6318c6318c6739ce7f53fffffff"),
                (x"ffffffffffa1ce318ce738c6318c6319ce739ce7f53fffffff"),
                (x"ffffffffffa0c6718ce739ce739ce739ce739ce7f53fffffff"),
                (x"ffffffffffa0c7e18ce739ce739ce739ce739fdef53fffffff"),
                (x"ffffffffffa1cfe18ce739ce739ce739ce739fdef53fffffff"),
                (x"ffffffffffa7bde38c7ef1ce739ce73fbc739fdef53fffffff"),
                (x"ffffffffffa7bde38c7ef1ce739ce73fbc739fdef53fffffff"),
                (x"ffffffffffa7bdef1c7ef1ce739ce7f7bc73fbdef53fffffff"),
                (x"fffffffffffd29ef1ce73f8e739ce7f1ce73fbdea53fffffff"),
                (x"fffffffffffd29ef78e73fbc739cfef1ce7f7bdea7ffffffff"),
                (x"ffffffffffffff4f7bc739e9ef7bd439cfef7a94ffffffffff"),
                (x"ffffffffffffff4f7bc739e9ef7bd439cfef7a94ffffffffff"),
                (x"fffffffffffffffa7bdef7a94a53d4f7bdef53ffffffffffff"),
                (x"fffffffffffffffa529defbb4a529405294a7a94ffffffffff"),
                (x"ffffffffffffff4f7a9defbde18fdef77bdf1fdea7ffffffff"),
                (x"ffffffffffffff43fa9defbdef7bdef7bd4f78e7f53fffffff"),
                (x"ffffffffffffff43fa9defbdef7bdef7bd4f78e7f53fffffff"),
                (x"fffffffffffd294f7a94a77def7a9ef77b4f53dea529ffffff"),
                (x"ffffffffffa529ea7a94a529def7b4a5294f53def529ffffff"),
                (x"ffffffffffa5294f7bc005294a5294a529e00294a53fffffff"),
                (x"ffffffffff0529da528005294ef7bda5294a53bda53fffffff"),
                (x"ffffffffff0529da528005294ef7bda5294a53bda53fffffff"),
                (x"fffffffffffd294ef694a78fea53c719cfe05294a7ffffffff"),
                (x"fffffffffff8014a5014a53d400014f7bd400000ffffffffff"),
                (x"fffffffffffffff00014a5294003c73d280fffffffffffffff"),
                (x"ffffffffffffffffffe005280f7a94f7bc0fffffffffffffff"),
                (x"ffffffffffffffffffe005280f7a94f7bc0fffffffffffffff"),
                (x"fffffffffffffffffffff8000f78e7a001ffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a529e07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a529407ffffffffffffffffff"),

                -- 3_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294f7bdef7bdffffffffffffffff"),
                (x"fffffffffffffffa53def1c6318c6339cfef7fffffffffffff"),
                (x"ffffffffffffff4f1ce739ce739c6318c633fbffffffffffff"),
                (x"fffffffffffd29e39ce739ce318c631fbcf1bfdeffffffffff"),
                (x"fffffffffffd29e39ce739ce318c631fbcf1bfdeffffffffff"),
                (x"fffffffffffd28739ce738c6318c63f0c63295efffffffffff"),
                (x"ffffffffffa7bc73f8e318cfef78fe1bdfe1d0a5a7ffffffff"),
                (x"ffffffffffa7bc7f78e73fbc7f7bc37fbc0180a5a7ffffffff"),
                (x"ffffffffffa7bc7f78e73fbc7f7bc37fbc0180a5a7ffffffff"),
                (x"fffffffff4f7bdef1cfef7a9418c7ef528078063a7ffffffff"),
                (x"fffffffff4f7bdef1fd4a51e37bfdef5280781efa7ffffffff"),
                (x"fffffffff4f7bdef780f7bfdef7bdef7bd4f51ef07ffffffff"),
                (x"fffffffff4f7bdef501ef7bdef7a800001ef7800ffffffffff"),
                (x"ffffffffffa7bdef7814a7bdea50190000000000ffffffffff"),
                (x"ffffffffffa7bdef7814a7bdea50190000000000ffffffffff"),
                (x"ffffffffffa7bdea7bd4a0294a5019ce72739c00ffffffffff"),
                (x"fffffffffffd29ea7a94a02947bc199ce6739c00ffffffffff"),
                (x"fffffffffffd294a5294a0294f79fe9d28329463ffffffffff"),
                (x"ffffffffffffffea5294a0294f7bcf18c6f780a5a7ffffffff"),
                (x"ffffffffffffffea5294a0294f7bcf18c6f780a5a7ffffffff"),
                (x"fffffffffffffffa5294a0294f7bdef3de078063a7ffffffff"),
                (x"fffffffffffffffffe94a5014a53def3df478000ffffffffff"),
                (x"ffffffffffffffff8294a528000014a5294003ffffffffffff"),
                (x"fffffffffffffff078f4a77d4a5294a001ffffffffffffffff"),
                (x"fffffffffffffff078f4a77d4a5294a001ffffffffffffffff"),
                (x"fffffffffffffffa1c7ef53beef7def529ffffffffffffffff"),
                (x"fffffffffffffe0f1fdef529eef7c73d280a7fffffffffffff"),
                (x"fffffffffffffe0a78e73fa94a53c73fbd4f53ffffffffffff"),
                (x"fffffffffffffe0a1fdded000a529ef5294f53ffffffffffff"),
                (x"fffffffffffffe0a1fdded000a529ef5294f53ffffffffffff"),
                (x"fffffffffffffff07bb4a53c7a529ded280a03ffffffffffff"),
                (x"fffffffffffffff05294a53de0029ef5280fffffffffffffff"),
                (x"ffffffffffffffff8294a529400294a529ffffffffffffffff"),
                (x"ffffffffffffffffd014a0000a528719cfffffffffffffffff"),
                (x"ffffffffffffffffd014a0000a528719cfffffffffffffffff"),
                (x"ffffffffffffffffd294a0014a50fef529ffffffffffffffff"),
                (x"ffffffffffffffff800007c00a53d4a5280fffffffffffffff"),
                (x"fffffffffffffffffffffffff003de39ce0fffffffffffffff"),

                -- 3_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffff98c6a5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffdef78e739ce7318d4a7fffffffffffff"),
                (x"fffffffffffffffa78e738c6318c6318c67f53ffffffffffff"),
                (x"ffffffffffffff4f1c6318c6318c6318c633fa94ffffffffff"),
                (x"ffffffffffffff4f1c6318c6318c6318c633fa94ffffffffff"),
                (x"fffffffffffd29e38c6319cfef7bc739ce319fdea7ffffffff"),
                (x"fffffffffffd28719ce73f9e5294aff7bde39fdea7ffffffff"),
                (x"ffffffffffa7bc339cef794a3a53c51bdfef7bdef53fffffff"),
                (x"ffffffffffa7bc339cef794a3a53c51bdfef7bdef53fffffff"),
                (x"ffffffffffa7bc3f1de52be83003d478c6ff7a94f53fffffff"),
                (x"ffffffffffa1cfe3bcaf78c03003c07fbc37fa94f53fffffff"),
                (x"ffffffffffa1cf4f15e318c03a53c07fbde1fa94a53fffffff"),
                (x"ffffffffffa000f7d3cf78e83a53d47fbdea3def053fffffff"),
                (x"ffffffffffa001ef001ef3c637bfcff7bc007bde053fffffff"),
                (x"ffffffffffa001ef001ef3c637bfcff7bc007bde053fffffff"),
                (x"ffffffffffa5294f032000294a52940001907a94a53fffffff"),
                (x"ffffffffffa5280a0339ce4e739ce7ce73905000a53fffffff"),
                (x"fffffffffff8000a53339cfd4a529e9ce79a500007ffffffff"),
                (x"fffffffffffffe0f53339f8a5294a3f4e79a7800ffffffffff"),
                (x"fffffffffffffe0f53339f8a5294a3f4e79a7800ffffffffff"),
                (x"fffffffffffffe0a7874a1463003cf1d28ff5000ffffffffff"),
                (x"fffffffffffd29ea79f4a3c03003c0f528ff53dea7ffffffff"),
                (x"ffffffffffa1ce7f53d4a3e83003d4f529ea7bdef7bdffffff"),
                (x"fffffffff4f1cfef7694a51eff7bdea529eefa94f1cfef7fff"),
                (x"fffffffff4f1cfef7694a51eff7bdea529eefa94f1cfef7fff"),
                (x"fffffffffe18c67f529ef7694a5294f77bea53de39c7ef53ff"),
                (x"ffffffd2833fbdda029ef50e739ce73d29e053dea53b4a53ff"),
                (x"ffffffd287ed294f5014a7bdef7bdef5294a5294a5294a7fff"),
                (x"fffffffff4a529e38e94a5294a5294a529407c00a7bd4a7fff"),
                (x"fffffffff4a529e38e94a5294a5294a529407c00a7bd4a7fff"),
                (x"ffffffffffa529e39e94a529def7b4a7bd407c00f1cf4a7fff"),
                (x"fffffffffff8014f5014a78e318cfef5294a7fffa78e007fff"),
                (x"fffffffffffffe000294a53c7f7a9419cfe07fff0001ffffff"),
                (x"fffffffffffffffffff4a5280a5067f7bd4fffffffffffffff"),
                (x"fffffffffffffffffff4a5280a5067f7bd4fffffffffffffff"),
                (x"ffffffffffffffffffe007a80a53def529ffffffffffffffff"),
                (x"fffffffffffffffffffff80000029ea001ffffffffffffffff"),
                (x"fffffffffffffffffffffffff000e307ffffffffffffffffff"),

                -- 3_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffdef7bdea5294a529ffffffffffffffff"),
                (x"ffffffffffffffff78e738c6318c67f7bd4a7fffffffffffff"),
                (x"ffffffffffffffe38c6318c6739ce739ce7f53ffffffffffff"),
                (x"ffffffffffffbcf1bfc318c6318ce739ce73fa94ffffffffff"),
                (x"ffffffffffffbcf1bfc318c6318ce739ce73fa94ffffffffff"),
                (x"fffffffffffbde528c7ef0c6318c6339ce739e94ffffffffff"),
                (x"ffffffffffa14b41f9e31f8fef78e319cfe39fdea7ffffffff"),
                (x"ffffffffffa14a0183cf78fde39fde39cfef1fdea7ffffffff"),
                (x"ffffffffffa14a0183cf78fde39fde39cfef1fdea7ffffffff"),
                (x"ffffffffffa0c607829ef7863a529ef1ce7f7bdef53fffffff"),
                (x"ffffffffffa3de07829ef7bcf18df4a7bc7f7bdef53fffffff"),
                (x"ffffffffff03df4f53def7bdef7bcf7801ef7bdef53fffffff"),
                (x"fffffffffff801ef78000029ef7bdef0014f7bdef53fffffff"),
                (x"fffffffffff80000000006414f7bdea001ef7bdea7ffffffff"),
                (x"fffffffffff80000000006414f7bdea001ef7bdea7ffffffff"),
                (x"fffffffffff800739f39ce414a5280a7bdea7bdea7ffffffff"),
                (x"fffffffffff800739e739e40fa5280a529ea7a94ffffffffff"),
                (x"fffffffffff8c6528e939f9fea5280a5294a5294ffffffffff"),
                (x"ffffffffffa14a07bc74a3fdea5280a5294a7bffffffffffff"),
                (x"ffffffffffa14a07bc74a3fdea5280a5294a7bffffffffffff"),
                (x"ffffffffffa0c60781f4a7bdea5280a5294a7fffffffffffff"),
                (x"fffffffffff80007d1f4a7bd4a5014a529ffffffffffffffff"),
                (x"fffffffffffffe005294a500000294a5280fffffffffffffff"),
                (x"fffffffffffffffffc14a5294a53dda1cfe07fffffffffffff"),
                (x"fffffffffffffffffc14a5294a53dda1cfe07fffffffffffff"),
                (x"fffffffffffffffffe9ef7bddf7bb4f0c67a7fffffffffffff"),
                (x"fffffffffffffffa028739fddf7a94f7bc7f03ffffffffffff"),
                (x"ffffffffffffff4f53c739fd4a529e39cfea03ffffffffffff"),
                (x"ffffffffffffff4f529ef7a9400014efbc7a03ffffffffffff"),
                (x"ffffffffffffff4f529ef7a9400014efbc7a03ffffffffffff"),
                (x"fffffffffffffe0a029def69439fd4a77be07fffffffffffff"),
                (x"ffffffffffffffff829ef7a80f7bd4a529407fffffffffffff"),
                (x"fffffffffffffffffe94a5280a5294a5280fffffffffffffff"),
                (x"fffffffffffffffffce319e9400000a0014fffffffffffffff"),
                (x"fffffffffffffffffce319e9400000a0014fffffffffffffff"),
                (x"fffffffffffffffffe9ef78f4a5000a5294fffffffffffffff"),
                (x"ffffffffffffffff8294a53d40001f00000fffffffffffffff"),
                (x"ffffffffffffffff80e73fbc0fffffffffffffffffffffffff"),

                -- 4_character_0_0
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c6318ca53ffffffffffff"),
                (x"fffffffffffd2946318c6318c6318c6319e63294a7ffffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"fffffffffffd2946318c6318c6318c6318c63294a7ffffffff"),
                (x"fffffffffffd2946318c6318c6318c6318c63294a7ffffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318c653fffffff"),
                (x"fffffffff4a31946318c6318c6318c6318c632946529ffffff"),
                (x"fffffffff4a31946318c6318c6318c6318c632946529ffffff"),
                (x"fffffffff4a528c633cc633cc6319ef318ca318ca529ffffff"),
                (x"fffffffff4a528ca318c633de6318c6318c6518ca529ffffff"),
                (x"fffffffff4a5294a318c6518c6318c6528c65294a529ffffff"),
                (x"fffffffff4a528ca5194a518c6328c6529465294a529ffffff"),
                (x"ffffffffff0528ca5194a528ca528ca5294a5294a03fffffff"),
                (x"ffffffffff0528ca5194a528ca528ca5294a5294a03fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294a03fffffff"),
                (x"fffffffffff8014a5194a5294a5294a5294a529407ffffffff"),
                (x"fffffffffffffe0a5194a5194a5194a5294a5000ffffffffff"),
                (x"fffffffffffffff0528c65194a5194a5294a03ffffffffffff"),
                (x"fffffffffffffff0528c65194a5194a5294a03ffffffffffff"),
                (x"ffffffffffffbcf20294a5294a5294a5294011eff7ffffffff"),
                (x"ffffffffff790810900005294a5294a00002042123ffffffff"),
                (x"ffffffffff2842109463182940029400c63e8421097fffffff"),
                (x"ffffffffef094a5253c31f86318c63f0c7ea10a5285fffffff"),
                (x"ffffffffef094a5253c31f86318c63f0c7ea10a5285fffffff"),
                (x"fffffffffe204212d3def0c6318c631fbdea1421093dffffff"),
                (x"ffffffffec4b18cf03a318c6318c6318c7d0798c6259ffffff"),
                (x"ffffffffe04dee9077ddefbc318c7ef77bee8129ba41ffffff"),
                (x"ffffffffff00000677bdefa94a5294f77bdeb000003fffffff"),
                (x"ffffffffff00000677bdefa94a5294f77bdeb000003fffffff"),
                (x"fffffffffffffff074e738c67ef4e319ce7e83ffffffffffff"),
                (x"fffffffffffffffff4e738c67ef4e319ce7effffffffffffff"),
                (x"fffffffffffffffff7a739cfdef7a739cfdeffffffffffffff"),
                (x"ffffffffffffffff83bdef7bd003bdef7bd07fffffffffffff"),
                (x"ffffffffffffffff83bdef7bd003bdef7bd07fffffffffffff"),
                (x"ffffffffffffffff83bde9fbd003bd3f7bd07fffffffffffff"),
                (x"fffffffffffffffffc0739ce0ffc0739ce0fffffffffffffff"),
                (x"fffffffffffffffffc1defba0ffc1df77a0fffffffffffffff"),

                -- 4_character_0_1
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c6318ca5294a7ffffffff"),
                (x"ffffffffffffff4a319ef318c6318c6318c6318c6529ffffff"),
                (x"fffffffffffd2946318c6318c631946318c63294a53fffffff"),
                (x"fffffffffffd28c6318c6798c63194a319ea318ca53fffffff"),
                (x"fffffffffffd28c6318c6798c63194a319ea318ca53fffffff"),
                (x"ffffffffffa528ca318c6328cf7a944d28ca518c653fffffff"),
                (x"ffffffffffa52946318c6328c63289ba53465294653fffffff"),
                (x"ffffffffffa528c6518c6328ca5137bdef74b294a53fffffff"),
                (x"ffffffffffa528c6518c6328ca5137bdef74b294a53fffffff"),
                (x"ffffffffffa3194a3194a328ca52f7bdef7ba694a53fffffff"),
                (x"ffffffffffa5294a3294a32944a58cf3197bdc00a7ffffffff"),
                (x"ffffffffff05294a5294a5294bdd8ca5294bdc00ffffffffff"),
                (x"ffffffffff05294a5294a5189bdd2500017bdc00ffffffffff"),
                (x"fffffffffffd294a52894d197bdd2400017bdc00ffffffffff"),
                (x"fffffffffffd294a52894d197bdd2400017bdc00ffffffffff"),
                (x"fffffffffff8014a52894d297bdee463197bdc00ffffffffff"),
                (x"fffffffffffffe0a5294a5297bdee4631976318ca7ffffffff"),
                (x"fffffffffffffff05294a5137bdeecbdeecf798c67ffffffff"),
                (x"ffffffffffffffff8294a5197bdef46319e63294ffffffffff"),
                (x"ffffffffffffffff8294a5197bdef46319e63294ffffffffff"),
                (x"fffffffffffffffffe94a528cbdef4a318c653ffffffffffff"),
                (x"ffffffffffffffffffc4210be6318ca5294a7fffffffffffff"),
                (x"fffffffffffffffff8810848fef6946001efffffffffffffff"),
                (x"ffffffffffffffff15e52bde5f78636319df7fffffffffffff"),
                (x"ffffffffffffffff15e52bde5f78636319df7fffffffffffff"),
                (x"ffffffffffffffff3c81084aff7bc365adef7fffffffffffff"),
                (x"ffffffffffffffff10bef798c0001eeb18cf7fffffffffffff"),
                (x"fffffffffffffff01597bdd37bdd201daccf7fffffffffffff"),
                (x"fffffffffffffff032f7bdef7bdee0f5accf7fffffffffffff"),
                (x"fffffffffffffff032f7bdef7bdee0f5accf7fffffffffffff"),
                (x"ffffffffffffffff8137bdd37bdd20edadefffffffffffffff"),
                (x"fffffffffffffffffc000318c000073f7bffffffffffffffff"),
                (x"fffffffffffffffffc1def7bdef4e7ef7bffffffffffffffff"),
                (x"ffffffffffffffffffe0077bd39c67efffffffffffffffffff"),
                (x"ffffffffffffffffffe0077bd39c67efffffffffffffffffff"),
                (x"ffffffffffffffffffe0077a718cfdffffffffffffffffffff"),
                (x"fffffffffffffffffffff83a318c60ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83be297c0ffffffffffffffffffff"),

                -- 4_character_0_2
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c65294a53ffffffffffff"),
                (x"fffffffffffd294633cc6318c6318c6318c65294a7ffffffff"),
                (x"ffffffffffa528c6319ef328c6318c6318cf318ca53fffffff"),
                (x"fffffffffffd2946318c6528cf799467bd463294a7ffffffff"),
                (x"fffffffffffd2946318c6528cf799467bd463294a7ffffffff"),
                (x"ffffffffffa528c65194a529463294a318ca318ca53fffffff"),
                (x"ffffffffffa318c65194a3134a528c4d28ca3294653fffffff"),
                (x"fffffffff4a31946528c65ee9a5197ba534a5294a329ffffff"),
                (x"fffffffff4a31946528c65ee9a5197ba534a5294a329ffffff"),
                (x"fffffffff46528ca2697bdef7632f7bdef44d294a529ffffff"),
                (x"fffffffff4a528ca5d37bdef7bdef7bdee9bd18ca529ffffff"),
                (x"fffffffff4a5294a319ef32f7bdef767bcc65294a529ffffff"),
                (x"fffffffff4a529463194a5297bdef4a528c63294a529ffffff"),
                (x"ffffffffff0253465ca0002f7bdef700005bb294483fffffff"),
                (x"ffffffffff0253465ca0002f7bdef700005bb294483fffffff"),
                (x"ffffffffff0253465c80002f7bdef700004bb294483fffffff"),
                (x"fffffffffff8014a5c8c632f7bdef763184bd29407ffffffff"),
                (x"fffffffffffffe0a5c8c6318cbdd8c63184bd000ffffffffff"),
                (x"fffffffffffbde5032f7bb3dea53de65ef7600a57fffffffff"),
                (x"fffffffffffbde5032f7bb3dea53de65ef7600a57fffffffff"),
                (x"ffffffffff790812d18c6798ca518cf318ca142123ffffffff"),
                (x"ffffffffef284212528c63194bde8c63194a1021095fffffff"),
                (x"ffffffbde4214af21694a528c63194a5294291ef2908f7ffff"),
                (x"fffff794bef1085797bef0c7ef7bc31fbdd2bca527bc52bfff"),
                (x"fffff794bef1085797bef0c7ef7bc31fbdd2bca527bc52bfff"),
                (x"fffff7b1894b184f03d4a0e8cb59941d29e078846252c63fff"),
                (x"fffff62537ba52c003c31d3a3633bda0c7e0018c4dee94b3ff"),
                (x"fffff625374def76028318c6cb598318c74032f7ba6e94b3ff"),
                (x"ffffff80094def7677d4a7bccb599ef529eeb2f7ba52007fff"),
                (x"ffffff80094def7677d4a7bccb599ef529eeb2f7ba52007fff"),
                (x"ffffffffe04def7074fef7bde633def7bc7e82f7ba41ffffff"),
                (x"ffffffffff00000ff4e738c6318c6319ce7efc00003fffffff"),
                (x"fffffffffffffffff7a738cfdef7a719cfdeffffffffffffff"),
                (x"ffffffffffffffff83a739cfd003a739cfd07fffffffffffff"),
                (x"ffffffffffffffff83a739cfd003a739cfd07fffffffffffff"),
                (x"ffffffffffffffff83a318cfd003a718c7d07fffffffffffff"),
                (x"fffffffffffffffffc1def7a0ffc1def7a0fffffffffffffff"),
                (x"ffffffffffffffffffbdefba0ffc1df77bdfffffffffffffff"),

                -- 4_character_0_3
                (x"fffffffffffffffa5294a318c63294a529ffffffffffffffff"),
                (x"fffffffffffffffa5294a318c63294a529ffffffffffffffff"),
                (x"ffffffffffa5294a318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf318ca53ffffffffffff"),
                (x"fffffffff4a528c6318c6518c6318c6318c65294ffffffffff"),
                (x"fffffffff4a318ca7994a518c6319e6318c63294ffffffffff"),
                (x"fffffffff4a318ca7994a518c6319e6318c63294ffffffffff"),
                (x"fffffffff463194a32894d29e6328c6318ca3294a7ffffffff"),
                (x"fffffffff46529465137ba68c6328c6318c65294a7ffffffff"),
                (x"fffffffff4a528c4def7bdd346328c6319463294a7ffffffff"),
                (x"fffffffff4a528c4def7bdd346328c6319463294a7ffffffff"),
                (x"fffffffff4a5289bdef7bdef46328ca318ca518ca7ffffffff"),
                (x"ffffffffffa0017bdd9ef3189a528ca528ca5294a7ffffffff"),
                (x"fffffffffff8017bd294a3197a5294a5294a529407ffffffff"),
                (x"fffffffffff8017bdc00015374a594a5294a529407ffffffff"),
                (x"fffffffffff8017bdc0001137bdd944d294a5000ffffffffff"),
                (x"fffffffffff8017bdc0001137bdd944d294a5000ffffffffff"),
                (x"fffffffffff8017bdd8c612f7bde944d294a5000ffffffffff"),
                (x"ffffffffffa318c65d8c612f7bde94a5294a03ffffffffffff"),
                (x"ffffffffff6319ef32f7bb2f7bdd34a529407fffffffffffff"),
                (x"ffffffffff6528c6798c652f7bdd94a5280fffffffffffffff"),
                (x"ffffffffff6528c6798c652f7bdd94a5280fffffffffffffff"),
                (x"fffffffffffd29463194a52f763294a529ffffffffffffffff"),
                (x"fffffffffffffffa5294a318cf78a427bdffffffffffffffff"),
                (x"fffffffffffffffff80c6529d7bc810909efffffffffffffff"),
                (x"ffffffffffffffff758c60c7e295ef2bde5f7fffffffffffff"),
                (x"ffffffffffffffff758c60c7e295ef2bde5f7fffffffffffff"),
                (x"ffffffffffffffff7acc60fde7bca10908ff7fffffffffffff"),
                (x"ffffffffffffffff319def8006319ef14a4f7fffffffffffff"),
                (x"ffffffffffffffff32c318137bdd37bb18507fffffffffffff"),
                (x"ffffffffffffffff32def02f7bdef7bdeec07fffffffffffff"),
                (x"ffffffffffffffff32def02f7bdef7bdeec07fffffffffffff"),
                (x"fffffffffffffffffadde8137bdd37ba520fffffffffffffff"),
                (x"ffffffffffffffffffa739c006318c0001ffffffffffffffff"),
                (x"ffffffffffffffffffbde9cfdef7bde801ffffffffffffffff"),
                (x"fffffffffffffffffffde9c67ef7bd07ffffffffffffffffff"),
                (x"fffffffffffffffffffde9c67ef7bd07ffffffffffffffffff"),
                (x"ffffffffffffffffffffff4e339fbd07ffffffffffffffffff"),
                (x"fffffffffffffffffffff806318fa0ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83c5f7ba0ffffffffffffffffffff"),

                -- 4_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c6318ca53ffffffffffff"),
                (x"fffffffffffd2946318c6318c6318c6319e63294a7ffffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"fffffffffffd2946318c6318c6318c6318c63294a7ffffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318c653fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318c653fffffff"),
                (x"fffffffff4a31946318c6318c6318c6318c632946529ffffff"),
                (x"fffffffff4a528c633cc633cc6319ef318ca318ca529ffffff"),
                (x"fffffffff4a528ca318c633de6318c6318c6518ca529ffffff"),
                (x"fffffffff4a5294a318c6518c6318c6528c65294a529ffffff"),
                (x"fffffffff4a528ca5194a518c6328c6529465294a529ffffff"),
                (x"fffffffff4a528ca5194a518c6328c6529465294a529ffffff"),
                (x"ffffffffff0528ca5194a528ca528ca5294a5294a03fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294a03fffffff"),
                (x"fffffffffff8014a5194a5294a5294a5294a529407ffffffff"),
                (x"fffffffffffffe0a5194a5194a5194a5294a5000ffffffffff"),
                (x"fffffffffffffe0a5194a5194a5194a5294a5000ffffffffff"),
                (x"ffffffffffffffe0528c65194a5194a5294a03ffffffffffff"),
                (x"ffffffffffffbc520294a5294a5294a5294013deffffffffff"),
                (x"fffffffffff14a42740005294a5294a000008484f7ffffffff"),
                (x"fffffffffff10852d063182940029407bdd08421f7ffffffff"),
                (x"fffffffffff10852d063182940029407bdd08421f7ffffffff"),
                (x"fffffffffff14a42787ef0c6318fc31fbdd084842fbfffffff"),
                (x"ffffffffff67bdef53c318c6318fdd1fbd42948427bfffffff"),
                (x"ffffffffff0318c053bef0c6318c7eef7b408421f33fffffff"),
                (x"fffffffffff800007a9def7deef7bef7bc0f7bde4b3fffffff"),
                (x"fffffffffff800007a9def7deef7bef7bc0f7bde4b3fffffff"),
                (x"fffffffffffffffff7bde9cfdef7bdef7bd6252907ffffffff"),
                (x"fffffffffffffffff7bde9c63ef7a73f7bde8000ffffffffff"),
                (x"fffffffffffffffff7bdef4e7ef7bdef7a007fffffffffffff"),
                (x"fffffffffffffffffc1def7bd39c1de801ffffffffffffffff"),
                (x"fffffffffffffffffc1def7bd39c1de801ffffffffffffffff"),
                (x"ffffffffffffffffffe0074e7ef40007ffffffffffffffffff"),
                (x"fffffffffffffffffffff83c3f781fffffffffffffffffffff"),
                (x"fffffffffffffffffffff83ddef41fffffffffffffffffffff"),

                -- 4_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c6318ca5294a7ffffffff"),
                (x"ffffffffffffff4a319ef318c6318c6318c6318c6529ffffff"),
                (x"fffffffffffd2946318c6318c631946318c63294a53fffffff"),
                (x"fffffffffffd2946318c6318c631946318c63294a53fffffff"),
                (x"fffffffffffd28c6318c6798c63194a319ea318ca53fffffff"),
                (x"ffffffffffa528ca318c6328cf7a944d28ca518c653fffffff"),
                (x"ffffffffffa52946318c6328c63289ba53465294653fffffff"),
                (x"ffffffffffa52946318c6328c63289ba53465294653fffffff"),
                (x"ffffffffffa528c6518c6328ca5137bdef74b294a53fffffff"),
                (x"ffffffffffa3194a3194a328ca52f7bdef7ba694a53fffffff"),
                (x"ffffffffffa5294a3294a32944a58cf3197bdc00a7ffffffff"),
                (x"ffffffffff05294a5294a5294bdd8ca5294bdc00ffffffffff"),
                (x"ffffffffff05294a5294a5189bdd2500017bdc00ffffffffff"),
                (x"ffffffffff05294a5294a5189bdd2500017bdc00ffffffffff"),
                (x"fffffffffffd294a52894d197bdd2400017bdc00ffffffffff"),
                (x"fffffffffff8014a52894d297bdee463197bdc00ffffffffff"),
                (x"fffffffffffffe0a5294a5297bdee4631976318ca7ffffffff"),
                (x"fffffffffffffff05294a5137bdeecbdeecf798c67ffffffff"),
                (x"fffffffffffffff05294a5137bdeecbdeecf798c67ffffffff"),
                (x"ffffffffffffffff8294a5197bdef46319e6329467ffffffff"),
                (x"fffffffffffffffffe94a528cbdef4a318c65294ffffffffff"),
                (x"ffffffffffffffff83c5290af6318ca5294a7fffffffffffff"),
                (x"ffffffffffffffff80a420425f7a94a001efffffffffffffff"),
                (x"ffffffffffffffff80a420425f7a94a001efffffffffffffff"),
                (x"fffffffffffffff07884214a4a53def7bcc07fffffffffffff"),
                (x"fffffffffffffff078af78421f7bbef7bcc07fffffffffffff"),
                (x"fffffffffffffff051e4215fef78000529d67fffffffffffff"),
                (x"fffffffffffffff053c52f989632f7b801d67fffffffffffff"),
                (x"fffffffffffffff053c52f989632f7b801d67fffffffffffff"),
                (x"fffffffffffffff07a80026f74a6f7b801467fffffffffffff"),
                (x"fffffffffffffffe83def01374a537677a0fffffffffffffff"),
                (x"fffffffffffffffef4e73f40c63000077bffffffffffffffff"),
                (x"fffffffffffffff074e319fbd003bdefffffffffffffffffff"),
                (x"fffffffffffffff074e319fbd003bdefffffffffffffffffff"),
                (x"fffffffffffffff077a73f7bd003a73f7bffffffffffffffff"),
                (x"ffffffffffffffff80e319fa00001df7bdffffffffffffffff"),
                (x"ffffffffffffffff83bef17c0fffffffffffffffffffffffff"),

                -- 4_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c65294a53ffffffffffff"),
                (x"fffffffffffd294633cc6318c6318c6318c65294a7ffffffff"),
                (x"ffffffffffa528c6319ef328c6318c6318cf318ca53fffffff"),
                (x"ffffffffffa528c6319ef328c6318c6318cf318ca53fffffff"),
                (x"fffffffffffd2946318c6528cf799467bd463294a7ffffffff"),
                (x"ffffffffffa528c65194a529463294a318ca318ca53fffffff"),
                (x"ffffffffffa318c65194a3134a528c4d28ca3294653fffffff"),
                (x"ffffffffffa318c65194a3134a528c4d28ca3294653fffffff"),
                (x"fffffffff4a31946528c65ee9a5197ba534a5294a329ffffff"),
                (x"fffffffff46528ca2697bdef7632f7bdef44d294a529ffffff"),
                (x"fffffffff4a528ca5d37bdef7bdef7bdee9bd18ca529ffffff"),
                (x"fffffffff4a5294a319ef32f7bdef767bcc65294a529ffffff"),
                (x"fffffffff4a529463194a5297bdef4a528c63294a529ffffff"),
                (x"fffffffff4a529463194a5297bdef4a528c63294a529ffffff"),
                (x"ffffffffff0253465ca0002f7bdef700005bb294483fffffff"),
                (x"ffffffffff0253465c80002f7bdef700004bb294483fffffff"),
                (x"fffffffffff8014a5c8c632f7bdef763184bd29407ffffffff"),
                (x"fffffffffffffe0a5c8c6318cbdd8c63184bd000ffffffffff"),
                (x"fffffffffffffe0a5c8c6318cbdd8c63184bd000ffffffffff"),
                (x"ffffffffffffbcf032f7bb3dea53de65ef7603def7ffffffff"),
                (x"ffffffffff794a42d18c6798ca518cf318ca142127bfffffff"),
                (x"ffffffffef290842528c63194bde8c63194a0484217dffffff"),
                (x"fffffffbc423de521294a528c63194a5294ebc21090bef7fff"),
                (x"fffffffbc423de521294a528c63194a5294ebc21090bef7fff"),
                (x"fffffffbcf2908f7f69ef0c7ef7bc31fbd4a11ef7bcbef7fff"),
                (x"ffffffb18963de5053d4a0e8cb59941d29ea01294b3dffffff"),
                (x"ffffffb1894b18c053c31d3a3633bda0c60032f7ba59ffffff"),
                (x"ffffffb197ba520fd3a318c6cb59831f7acbdef74a59ffffff"),
                (x"ffffffb197ba520fd3a318c6cb59831f7acbdef74a59ffffff"),
                (x"ffffffb189bb180ff7def77ccb599df7bccbdd296301ffffff"),
                (x"ffffff80094b19fff4e738c63630e73f7a04dd8c003fffffff"),
                (x"ffffffffe00001fff7a738c67ef7bdef7bd00000ffffffffff"),
                (x"ffffffffffffffffffa739c6739c1def7bdfffffffffffffff"),
                (x"ffffffffffffffffffa739c6739c1def7bdfffffffffffffff"),
                (x"fffffffffffffffffffde8c6339c1def7bffffffffffffffff"),
                (x"ffffffffffffffffffe0077bdef40007ffffffffffffffffff"),
                (x"ffffffffffffffffffffff7beef7ffffffffffffffffffffff"),

                -- 4_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa5294a318c63294a529ffffffffffffffff"),
                (x"ffffffffffa5294a318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf318ca53ffffffffffff"),
                (x"fffffffff4a528c6318c6518c6318c6318c65294ffffffffff"),
                (x"fffffffff4a528c6318c6518c6318c6318c65294ffffffffff"),
                (x"fffffffff4a318ca7994a518c6319e6318c63294ffffffffff"),
                (x"fffffffff463194a32894d29e6328c6318ca3294a7ffffffff"),
                (x"fffffffff46529465137ba68c6328c6318c65294a7ffffffff"),
                (x"fffffffff46529465137ba68c6328c6318c65294a7ffffffff"),
                (x"fffffffff4a528c4def7bdd346328c6319463294a7ffffffff"),
                (x"fffffffff4a5289bdef7bdef46328ca318ca518ca7ffffffff"),
                (x"ffffffffffa0017bdd9ef3189a528ca528ca5294a7ffffffff"),
                (x"fffffffffff8017bd294a3197a5294a5294a529407ffffffff"),
                (x"fffffffffff8017bdc00015374a594a5294a529407ffffffff"),
                (x"fffffffffff8017bdc00015374a594a5294a529407ffffffff"),
                (x"fffffffffff8017bdc0001137bdd944d294a5000ffffffffff"),
                (x"fffffffffff8017bdd8c612f7bde944d294a5000ffffffffff"),
                (x"ffffffffffa318c65d8c612f7bde94a5294a03ffffffffffff"),
                (x"ffffffffff6319ef32f7bb2f7bdd34a529407fffffffffffff"),
                (x"ffffffffff6319ef32f7bb2f7bdd34a529407fffffffffffff"),
                (x"ffffffffff6528c6798c652f7bdd94a5280fffffffffffffff"),
                (x"fffffffffffd29463194a52f763294a529ffffffffffffffff"),
                (x"fffffffffffffffa5294a318c7bca42fbc0fffffffffffffff"),
                (x"fffffffffffffffff814a529e29421214a0fffffffffffffff"),
                (x"fffffffffffffffff814a529e29421214a0fffffffffffffff"),
                (x"fffffffffffffff033def7bd4210a52109e07fffffffffffff"),
                (x"fffffffffffffff033def7bbe08421794be07fffffffffffff"),
                (x"fffffffffffffff676800001ef79e523df407fffffffffffff"),
                (x"fffffffffffffff67417bdeec4a59e2fbd407fffffffffffff"),
                (x"fffffffffffffff67417bdeec4a59e2fbd407fffffffffffff"),
                (x"fffffffffffffff65017bdee9bdee903dfe07fffffffffffff"),
                (x"ffffffffffffffff83ac65d29bdd20f7bc0effffffffffffff"),
                (x"ffffffffffffffffffa00000c6301d39cfdeffffffffffffff"),
                (x"fffffffffffffffffffdef7a0ef7a719cfd07fffffffffffff"),
                (x"fffffffffffffffffffdef7a0ef7a719cfd07fffffffffffff"),
                (x"ffffffffffffffffffa739fa0ef7bd3f7bd07fffffffffffff"),
                (x"ffffffffffffffffffdef7400003a719ce0fffffffffffffff"),
                (x"fffffffffffffffffffffffff003c5f77a0fffffffffffffff"),

                -- 4_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c6318ca53ffffffffffff"),
                (x"fffffffffffd2946318c6318c6318c6319e63294a7ffffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"fffffffffffd2946318c6318c6318c6318c63294a7ffffffff"),
                (x"ffffffffffa528c6318c6318c6318c6318c6318ca53fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318c653fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318c653fffffff"),
                (x"fffffffff4a31946318c6318c6318c6318c632946529ffffff"),
                (x"fffffffff4a528c633cc633cc6319ef318ca318ca529ffffff"),
                (x"fffffffff4a528ca318c633de6318c6318c6518ca529ffffff"),
                (x"fffffffff4a5294a318c6518c6318c6528c65294a529ffffff"),
                (x"fffffffff4a528ca5194a518c6328c6529465294a529ffffff"),
                (x"fffffffff4a528ca5194a518c6328c6529465294a529ffffff"),
                (x"ffffffffff0528ca5194a528ca528ca5294a5294a03fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294a03fffffff"),
                (x"fffffffffff8014a5194a5294a5294a5294a529407ffffffff"),
                (x"fffffffffffffe0a5194a5194a5194a5294a5000ffffffffff"),
                (x"fffffffffffffe0a5194a5194a5194a5294a5000ffffffffff"),
                (x"fffffffffffffff0528c65194a5194a5294a03deffffffffff"),
                (x"ffffffffffffffe20294a5294a5294a5294013bdf7ffffffff"),
                (x"ffffffffffffbc40840005294a5294a0000e9084efbfffffff"),
                (x"ffffffffffffbc1087bef02940029400c63a14a527bfffffff"),
                (x"ffffffffffffbc1087bef02940029400c63a14a527bfffffff"),
                (x"fffffffffff14a4087bef0c7e18c631fbc3f10842fbfffffff"),
                (x"fffffffffff10842969ef0fbe18c6318c7ea7bdef33fffffff"),
                (x"ffffffffff67bc10869def7c318c631fbdda018c603fffffff"),
                (x"ffffffffff6253ef781ef7bddef7deef7b4f000007ffffffff"),
                (x"ffffffffff6253ef781ef7bddef7deef7b4f000007ffffffff"),
                (x"fffffffffff80094b3bdef7bdef7a73f7bdeffffffffffffff"),
                (x"fffffffffffffe0077bde9cfdef4633f7bdeffffffffffffff"),
                (x"ffffffffffffffff801def7bdef4e7ef7bdeffffffffffffff"),
                (x"ffffffffffffffffffe0077a039fbdef7a0fffffffffffffff"),
                (x"ffffffffffffffffffe0077a039fbdef7a0fffffffffffffff"),
                (x"fffffffffffffffffffff8000ef4e7e801ffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f787e07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0ef7be07ffffffffffffffffff"),

                -- 4_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c6318ca5294a7ffffffff"),
                (x"ffffffffffffff4a319ef318c6318c6318c6318c6529ffffff"),
                (x"fffffffffffd2946318c6318c631946318c63294a53fffffff"),
                (x"fffffffffffd2946318c6318c631946318c63294a53fffffff"),
                (x"fffffffffffd28c6318c6798c63194a319ea318ca53fffffff"),
                (x"ffffffffffa528ca318c6328cf7a944d28ca518c653fffffff"),
                (x"ffffffffffa52946318c6328c63289ba53465294653fffffff"),
                (x"ffffffffffa52946318c6328c63289ba53465294653fffffff"),
                (x"ffffffffffa528c6518c6328ca5137bdef74b294a53fffffff"),
                (x"ffffffffffa3194a3194a328ca52f7bdef7ba694a53fffffff"),
                (x"ffffffffffa5294a3294a32944a58cf3197bdc00a7ffffffff"),
                (x"ffffffffff05294a5294a5294bdd8ca5294bdc00ffffffffff"),
                (x"ffffffffff05294a5294a5189bdd2500017bdc00ffffffffff"),
                (x"ffffffffff05294a5294a5189bdd2500017bdc00ffffffffff"),
                (x"fffffffffffd294a52894d197bdd2400017bdc00ffffffffff"),
                (x"fffffffffff8014a52894d297bdee463197bdc00ffffffffff"),
                (x"fffffffffffffe0a5294a5297bdee4631976318ca7ffffffff"),
                (x"fffffffffffffff05294a5137bdeecbdeecf798c67ffffffff"),
                (x"fffffffffffffff05294a5137bdeecbdeecf798c67ffffffff"),
                (x"ffffffffffffffff8294a5197bdef46319e6329467ffffffff"),
                (x"fffffffffffffffffe94a528cbdef4a318c65294ffffffffff"),
                (x"ffffffffffffffff80a4217de6318ca5294a7fffffffffffff"),
                (x"fffffffffffffff01421091fdf7a944801efffffffffffffff"),
                (x"fffffffffffffff01421091fdf7a944801efffffffffffffff"),
                (x"ffffffffffffffff3c84207be18c7e67bddf7fffffffffffff"),
                (x"fffffffffffffe079021097bda506cb7bdd67fffffffffffff"),
                (x"fffffffffffffe02f9ef793d4f7bcc677be4b3ffffffffffff"),
                (x"fffffffffffffe0f26f7ba400f7bccb77be483ffffffffffff"),
                (x"fffffffffffffe0f26f7ba400f7bccb77be483ffffffffffff"),
                (x"fffffffffffffff026f7bdee9f7bacb7bc007fffffffffffff"),
                (x"fffffffffffffff03137bdef7000ecb77a0fffffffffffffff"),
                (x"ffffffffffffffff800c626e900063677bffffffffffffffff"),
                (x"ffffffffffffffff83bde8000ef4fdef7bffffffffffffffff"),
                (x"ffffffffffffffff83bde8000ef4fdef7bffffffffffffffff"),
                (x"fffffffffffffffff7bde8000ef4e319cfffffffffffffffff"),
                (x"ffffffffffffffff801def400003a7ef7a0fffffffffffffff"),
                (x"fffffffffffffffffffffffff003be2fbc0fffffffffffffff"),

                -- 4_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a5294fffffffffffffff"),
                (x"fffffffffffffffa528c6318c6318c65294a53ffffffffffff"),
                (x"fffffffffffd294633cc6318c6318c6318c65294a7ffffffff"),
                (x"ffffffffffa528c6319ef328c6318c6318cf318ca53fffffff"),
                (x"ffffffffffa528c6319ef328c6318c6318cf318ca53fffffff"),
                (x"fffffffffffd2946318c6528cf799467bd463294a7ffffffff"),
                (x"ffffffffffa528c65194a529463294a318ca318ca53fffffff"),
                (x"ffffffffffa318c65194a3134a528c4d28ca3294653fffffff"),
                (x"ffffffffffa318c65194a3134a528c4d28ca3294653fffffff"),
                (x"fffffffff4a31946528c65ee9a5197ba534a5294a329ffffff"),
                (x"fffffffff46528ca2697bdef7632f7bdef44d294a529ffffff"),
                (x"fffffffff4a528ca5d37bdef7bdef7bdee9bd18ca529ffffff"),
                (x"fffffffff4a5294a319ef32f7bdef767bcc65294a529ffffff"),
                (x"fffffffff4a529463194a5297bdef4a528c63294a529ffffff"),
                (x"fffffffff4a529463194a5297bdef4a528c63294a529ffffff"),
                (x"ffffffffff0253465ca0002f7bdef700005bb294483fffffff"),
                (x"ffffffffff0253465c80002f7bdef700004bb294483fffffff"),
                (x"fffffffffff8014a5c8c632f7bdef763184bd29407ffffffff"),
                (x"fffffffffffffe0a5c8c6318cbdd8c63184bd000ffffffffff"),
                (x"fffffffffffffe0a5c8c6318cbdd8c63184bd000ffffffffff"),
                (x"ffffffffffffbde032f7bb3dea53de65ef7601eff7ffffffff"),
                (x"fffffffffff10812d18c6798ca518cf318ca14842bffffffff"),
                (x"fffffffffe290840d28c63194bde8c63194a1084215fffffff"),
                (x"fffffffbc52042179694a528c63194a5294f10a57909ef7fff"),
                (x"fffffffbc52042179694a528c63194a5294f10a57909ef7fff"),
                (x"fffffffbc57bdef2529ef0c7ef7bc31fbd4ed1ef215fef7fff"),
                (x"fffffffffe62529053d4a0e8cb59941d29ea00a57b12c67fff"),
                (x"ffffffffec4def7600031d3a3633bda0c7ea018c6252c67fff"),
                (x"ffffffffec4a537bdd9de8c6cb598318c7da7c004deec67fff"),
                (x"ffffffffec4a537bdd9de8c6cb598318c7da7c004deec67fff"),
                (x"ffffffffe063189bdd9ef7bacb599eefbdeefc0065d2c67fff"),
                (x"ffffffffff0000cba41de9ce3630e319ce7effff6252007fff"),
                (x"fffffffffffffe0003bdef7bdef4e319cfdeffff0001ffffff"),
                (x"ffffffffffffffffffbdef7a039ce339cfdfffffffffffffff"),
                (x"ffffffffffffffffffbdef7a039ce339cfdfffffffffffffff"),
                (x"fffffffffffffffffffdef7a039c631f7bffffffffffffffff"),
                (x"fffffffffffffffffffff8000ef7bde801ffffffffffffffff"),
                (x"fffffffffffffffffffffffffef7ddefffffffffffffffffff"),

                -- 4_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa5294a318c63294a529ffffffffffffffff"),
                (x"ffffffffffa5294a318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf318ca53ffffffffffff"),
                (x"fffffffff4a528c6318c6518c6318c6318c65294ffffffffff"),
                (x"fffffffff4a528c6318c6518c6318c6318c65294ffffffffff"),
                (x"fffffffff4a318ca7994a518c6319e6318c63294ffffffffff"),
                (x"fffffffff463194a32894d29e6328c6318ca3294a7ffffffff"),
                (x"fffffffff46529465137ba68c6328c6318c65294a7ffffffff"),
                (x"fffffffff46529465137ba68c6328c6318c65294a7ffffffff"),
                (x"fffffffff4a528c4def7bdd346328c6319463294a7ffffffff"),
                (x"fffffffff4a5289bdef7bdef46328ca318ca518ca7ffffffff"),
                (x"ffffffffffa0017bdd9ef3189a528ca528ca5294a7ffffffff"),
                (x"fffffffffff8017bd294a3197a5294a5294a529407ffffffff"),
                (x"fffffffffff8017bdc00015374a594a5294a529407ffffffff"),
                (x"fffffffffff8017bdc00015374a594a5294a529407ffffffff"),
                (x"fffffffffff8017bdc0001137bdd944d294a5000ffffffffff"),
                (x"fffffffffff8017bdd8c612f7bde944d294a5000ffffffffff"),
                (x"ffffffffffa318c65d8c612f7bde94a5294a03ffffffffffff"),
                (x"ffffffffff6319ef32f7bb2f7bdd34a529407fffffffffffff"),
                (x"ffffffffff6319ef32f7bb2f7bdd34a529407fffffffffffff"),
                (x"ffffffffff6528c6798c652f7bdd94a5280fffffffffffffff"),
                (x"fffffffffffd29463194a52f763294a529ffffffffffffffff"),
                (x"fffffffffffffffa5294a318cf7bc5214a0fffffffffffffff"),
                (x"fffffffffffffffff8094d29eef6840842507fffffffffffff"),
                (x"fffffffffffffffff8094d29eef6840842507fffffffffffff"),
                (x"ffffffffffffffff77cc67863f78a12108ff7fffffffffffff"),
                (x"fffffffffffffff677d6b3074ef4a508424783ffffffffffff"),
                (x"fffffffffffffec4fbac633dea53c47bdfe283ffffffffffff"),
                (x"fffffffffffffe04fbb6b33de00009bdee9f03ffffffffffff"),
                (x"fffffffffffffe04fbb6b33de00009bdee9f03ffffffffffff"),
                (x"fffffffffffffff003d6b33be4a6f7bdee907fffffffffffff"),
                (x"ffffffffffffffff83b6b30e0bdef7ba52c07fffffffffffff"),
                (x"ffffffffffffffffffac60c604a6e960000fffffffffffffff"),
                (x"ffffffffffffffffffbdef4fd00000ef7a0fffffffffffffff"),
                (x"ffffffffffffffffffbdef4fd00000ef7a0fffffffffffffff"),
                (x"fffffffffffffffffce318cfd00000ef7bdfffffffffffffff"),
                (x"ffffffffffffffff83bde9fa00001de8000fffffffffffffff"),
                (x"ffffffffffffffff83c52fba0fffffffffffffffffffffffff"),

                -- 5_character_0_0
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffff4ef5ce739ce739ce739ceef694ffffffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b9cd739ceed3fffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad6b5ae6b9ce7769ffffff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad739ce73bb4a7fff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad739ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad735ce739d4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4a7fff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad735ce6bbb4a7fff"),
                (x"ffffffd29deb9ce6b5ad6b5ad6b5ad6b5ad6b9ad777b4a7fff"),
                (x"ffffffd294ef7bd739cd6b5ad6b5ad6b5ad73bbdef694a7fff"),
                (x"fffffffff4ef7bdef7ae739ce739ce739ddef7bdef69ffffff"),
                (x"ffffffffffa529def7bdef7bdef7bdef7bdef7bded3bffffff"),
                (x"ffffffffffa529def7bdef7bdef7bdef7bdef7bded3bffffff"),
                (x"ffffffffffef7b4a53bdef7bdef7bdef7bda5294efffffffff"),
                (x"ffffffffffff7bda5294a53bdef7bda5294a529407ffffffff"),
                (x"fffffffffffffe0a77b4a77bdef7bded29ded000ffffffffff"),
                (x"fffffffffffffff053bdef7bdef7bded294a03ffffffffffff"),
                (x"fffffffffffffff053bdef7bdef7bded294a03ffffffffffff"),
                (x"ffffffffffffff4a529ded3b4ef69da5294a5294ffffffffff"),
                (x"fffffffffffd29da77b4a5294a5294a529ded3bda7ffffffff"),
                (x"ffffffffffa77beef7def7414a5280efbdeef7deed3fffffff"),
                (x"ffffffffff07bdef53def7bdef7bdef7bdea7bdef03fffffff"),
                (x"ffffffffff07bdef53def7bdef7bdef7bdea7bdef03fffffff"),
                (x"ffffffffec48014ed3bef7bd30867ef7bdda76940259ffffff"),
                (x"ffffffffec4dee0053bef7bdef7bdef7bdda0000ba59ffffff"),
                (x"ffffffffe04dee90529def7c19cc3eef7b4a0129ba41ffffff"),
                (x"ffffffffff00000a53b4a529da53b4a529da5000003fffffff"),
                (x"ffffffffff00000a53b4a529da53b4a529da5000003fffffff"),
                (x"fffffffffffffffa53bef7bdef7bdef7bdda53ffffffffffff"),
                (x"ffffffffffffffffd29defbdef7bdef77b4a7fffffffffffff"),
                (x"fffffffffffffffff3bdef7bde73bdef7bde7fffffffffffff"),
                (x"ffffffffffffffff83ae739dd003ae739dd07fffffffffffff"),
                (x"ffffffffffffffff83ae739dd003ae739dd07fffffffffffff"),
                (x"ffffffffffffffff838e73bbc0039d739dc07fffffffffffff"),
                (x"fffffffffffffffffc1ce77a0ffc1def380fffffffffffffff"),
                (x"fffffffffffffffffc0000000ffc0000000fffffffffffffff"),

                -- 5_character_0_1
                (x"ffffffffffffffffffffffe94ef7bdef7bdef7ffffffffffff"),
                (x"ffffffffffffffffffffffe94ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffe94a77ae739ad6b5ad73bbda7ffffffff"),
                (x"fffffffffffffffa77ae735ad6b5ad6b5ad6b5ceed3fffffff"),
                (x"fffffffffffd29deb9ad6b5ad6b5ad6b5ad6b5ad753fffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b5ad777bda53fffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b5ad777bda53fffffff"),
                (x"fffffffff4eb9ce6b9ad6b5ad6b5ae777bdefbbdeb3fffffff"),
                (x"fffffffff4739ce735cd6b5ae73bbded29def5291f7fffffff"),
                (x"ffffffd29d739ce739ae739ddef69df77bdedef767ffffffff"),
                (x"ffffffd29d739ce739ae739ddef69df77bdedef767ffffffff"),
                (x"ffffffd29d739ce739ce777b4ef7deef7b7bdd2907ffffffff"),
                (x"ffffffd29deb9ce73bb4a53bdef7bdbdef7bdd8c67ffffffff"),
                (x"ffffff8014a77bda53bded3bdbdd2c63197bdd8cffffffffff"),
                (x"ffffffffe0f5294a53bdef477bdd2500017bdc00ffffffffff"),
                (x"ffffffffffa77bded28948d37bdd2400017bdc00ffffffffff"),
                (x"ffffffffffa77bded28948d37bdd2400017bdc00ffffffffff"),
                (x"ffffffffffa319da5297b8d37bdee4ef7b7bdc00ffffffffff"),
                (x"ffffffffffa77b4ef694a3137bdee4f7bd7bdc00ffffffffff"),
                (x"fffffffffffd294eb3b4a5137bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffffffffa7694a5189bdef7bdef7ba400ffffffffff"),
                (x"fffffffffffffffa7694a5189bdef7bdef7ba400ffffffffff"),
                (x"ffffffffffffffffd294a528c4a6f7bdef7483ffffffffffff"),
                (x"fffffffffffffffff7bef77b46318c6318007fffffffffffff"),
                (x"fffffffffffffffef7def7a9def6800001ffffffffffffffff"),
                (x"fffffffffffffffefbdef7a9df7bb4a529dfffffffffffffff"),
                (x"fffffffffffffffefbdef7a9df7bb4a529dfffffffffffffff"),
                (x"fffffffffffffffed0b4a03b4f7bd4ed29dfffffffffffffff"),
                (x"fffffffffffffff0312c60294ef7a06d280fffffffffffffff"),
                (x"fffffffffffffff05ef7bb3debdee068000fffffffffffffff"),
                (x"fffffffffffffff026f7ba7debdee0a0000fffffffffffffff"),
                (x"fffffffffffffff026f7ba7debdee0a0000fffffffffffffff"),
                (x"fffffffffffffffef537ba694bdd3def7a0fffffffffffffff"),
                (x"fffffffffffffffed3a00529400014e001dfffffffffffffff"),
                (x"fffffffffffffffed29defbddef694e77a0fffffffffffffff"),
                (x"fffffffffffffff0529defbdda529de77a0fffffffffffffff"),
                (x"fffffffffffffff0529defbdda529de77a0fffffffffffffff"),
                (x"ffffffffffffffff801ce77ae739dde7ffffffffffffffffff"),
                (x"ffffffffffffffffffe00039def780ffffffffffffffffffff"),
                (x"fffffffffffffffffffff8014a5000ffffffffffffffffffff"),

                -- 5_character_0_2
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffff4eb9cd6b5ad6b5ad6b9dded294ffffffffff"),
                (x"ffffffffffa77ae6b5ad6b5ad6b5ad739ce777bded3fffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ae777ae73bbdef69ffffff"),
                (x"ffffffd29d739ce777bdefbdef7bdeed294a77bdef7b4a7fff"),
                (x"ffffffd29d739ce777bdefbdef7bdeed294a77bdef7b4a7fff"),
                (x"ffffffd29d739d4a77b4a77bdef7bded294a5294ef7b4a7fff"),
                (x"ffffffd294ef7bda77bdef58318d8cef7bded294ef7b4a7fff"),
                (x"ffffff8014ed29deb19dea58318c6c4f7acef7bda768007fff"),
                (x"ffffff8014ed29deb19dea58318c6c4f7acef7bda768007fff"),
                (x"ffffffffe0ef7bdea6f7bdee918d37bdef7677bdef41ffffff"),
                (x"fffffffff403183edef7bdef7bdef7bdef7bf463e829ffffff"),
                (x"fffffffff460c6ceb2f7bdef7bdef7bdef76758c1f69ffffff"),
                (x"ffffffffffeb19d4a6f7bdef7bdef7bdef74a694677fffffff"),
                (x"ffffffffffa319d4dd8c632f7bdef76318c4a694653fffffff"),
                (x"ffffffffffa319d4dd8c632f7bdef76318c4a694653fffffff"),
                (x"ffffffffff0529d4dca0002f7bdef700005ba694a03fffffff"),
                (x"ffffffffff05ef44dc80002f7bdef700004ba694b83fffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"ffffffffffffffd026f7bdef7bdef7bdef7483bdffffffffff"),
                (x"ffffffffffed29da3137bdef7bdef7bdee9653bda77fffffff"),
                (x"fffffffffdefbdded3ac62537bdee94b19da77bdf77bffffff"),
                (x"fffffff7bdf7bdda53bded18c6318ca77bda53bdf7bbdeffff"),
                (x"fffffff7bdf7bdda53bded18c6318ca77bda53bdf7bbdeffff"),
                (x"ffffff8000a5294a53bef7a80a5014f7bdda5294a500007fff"),
                (x"fffff62537bb194ed3def7bada51bdf7bdea769465ee94b3ff"),
                (x"fffff6252cf5294053bef780def5a0f7bdda0294a79894b3ff"),
                (x"ffffff801ea252c0769def81400280f77b4e818c4d3c007fff"),
                (x"ffffff801ea252c0769def81400280f77b4e818c4d3c007fff"),
                (x"ffffff8014bdee965294a53bdef7bda5294a3129bde8007fff"),
                (x"ffffffffe0bdee9053bdef414ef680ef7bda0129bdc1ffffff"),
                (x"ffffffffff00000053bef781d73ba0f7bdda0000003fffffff"),
                (x"fffffffffffffffff7bdef5dce738eef7bdeffffffffffffff"),
                (x"fffffffffffffffff7bdef5dce738eef7bdeffffffffffffff"),
                (x"fffffffffffffffff3ad6b5dd003ae6b5bde7fffffffffffff"),
                (x"ffffffffffffffff83ae73bbd003bd739dd07fffffffffffff"),
                (x"fffffffffffffffffe94a5294ffe94a5294fffffffffffffff"),

                -- 5_character_0_3
                (x"ffffffffffffffdef7bdef7bda529fffffffffffffffffffff"),
                (x"ffffffffffffffdef7bdef7bda529fffffffffffffffffffff"),
                (x"ffffffffffa77ae735ad6b5ae73bbda529ffffffffffffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad777bda77ffffffffffff"),
                (x"fffffffff4735ad6b5ad6b5ad6b5ad6b5aeef694ffffffffff"),
                (x"fffffffff4a77bd735ad6b5ad6b5ad6b5ad73bbda7ffffffff"),
                (x"fffffffff4a77bd735ad6b5ad6b5ad6b5ad73bbda7ffffffff"),
                (x"ffffffffecef7beef7ae739ad6b5ad6b5ae6b9ceed3fffffff"),
                (x"fffffffffd1a53def69def7ae739ad6b9cd739ce753fffffff"),
                (x"ffffffffff65ef7ef7bef769def5ce735ae739ce7769ffffff"),
                (x"ffffffffff65ef7ef7bef769def5ce735ae739ce7769ffffff"),
                (x"ffffffffff02537bdfbdef7dda53bd739ce739ce7769ffffff"),
                (x"ffffffffff63197bdef7bdfbdef7b4a77ae739ceef69ffffff"),
                (x"fffffffffffb197bdd8c63137ef7b4ef7b4a77bda501ffffff"),
                (x"fffffffffff8017bdc0001537bdc63677b4a5294f03fffffff"),
                (x"fffffffffff8017bdc0001137bdd234d294ef7bda7ffffffff"),
                (x"fffffffffff8017bdc0001137bdd234d294ef7bda7ffffffff"),
                (x"fffffffffff8017bdfbde92f7bdd23bd294a758ca7ffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd2ca529ded3bda7ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a77aced294ffffffffff"),
                (x"fffffffffff8009bdef7bdef74a594a529da7fffffffffffff"),
                (x"fffffffffff8009bdef7bdef74a594a529da7fffffffffffff"),
                (x"fffffffffffffe04def7bdee963294a5294fffffffffffffff"),
                (x"fffffffffffffff0018c6318ca53bdf77bdfffffffffffffff"),
                (x"fffffffffffffffffc000029def69ef7bddeffffffffffffff"),
                (x"fffffffffffffffff694a53beef69ef7bdeeffffffffffffff"),
                (x"fffffffffffffffff694a53beef69ef7bdeeffffffffffffff"),
                (x"fffffffffffffffff69ded3dea53a0a77b4effffffffffffff"),
                (x"ffffffffffffffff828d683bda52806252c07fffffffffffff"),
                (x"ffffffffffffffff800d682f7f7bccbdef707fffffffffffff"),
                (x"ffffffffffffffff8014a02f7f7bc9bdee907fffffffffffff"),
                (x"ffffffffffffffff8014a02f7f7bc9bdee907fffffffffffff"),
                (x"ffffffffffffffff83bdef537a5289ba53deffffffffffffff"),
                (x"fffffffffffffffff41ce5000a5294077b4effffffffffffff"),
                (x"ffffffffffffffff83bce529def7deed294effffffffffffff"),
                (x"ffffffffffffffff83bce7694ef7deed29407fffffffffffff"),
                (x"ffffffffffffffff83bce7694ef7deed29407fffffffffffff"),
                (x"fffffffffffffffffffce75ce73bbde0000fffffffffffffff"),
                (x"fffffffffffffffffffff839def78007ffffffffffffffffff"),
                (x"fffffffffffffffffffff8014a5000ffffffffffffffffffff"),

                -- 5_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffff4ef5ce739ce739ce739ceef694ffffffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b9cd739ceed3fffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b9cd739ceed3fffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad6b5ae6b9ce7769ffffff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad739ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad735ce739d4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4a7fff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad735ce6bbb4a7fff"),
                (x"ffffffd29deb9ce6b5ad6b5ad6b5ad6b5ad6b9ad777b4a7fff"),
                (x"ffffffd294ef7bd739cd6b5ad6b5ad6b5ad73bbdef694a7fff"),
                (x"ffffffd294ef7bd739cd6b5ad6b5ad6b5ad73bbdef694a7fff"),
                (x"fffffffff4ef7bdef7ae739ce739ce739ddef7bdef69ffffff"),
                (x"ffffffffffa529def7bdef7bdef7bdef7bdef7bded3bffffff"),
                (x"ffffffffffef7b4a53bdef7bdef7bdef7bda5294ef7fffffff"),
                (x"ffffffffffff7bda5294a53bdef7bda5294a53bd07ffffffff"),
                (x"ffffffffffff7bda5294a53bdef7bda5294a53bd07ffffffff"),
                (x"fffffffffffffe0ef7b4a77bdef7bded29def400ffffffffff"),
                (x"fffffffffffffff053ac65194ef7bdef7aca03ffffffffffff"),
                (x"fffffffffffd294ed29ded3b4ef69da5294a5294ffffffffff"),
                (x"ffffffffffa529ef7694a5294a52940529df7a94a7ffffffff"),
                (x"ffffffffffa529ef7694a5294a52940529df7a94a7ffffffff"),
                (x"ffffffffff07bdef53bef7694a5280a529df7bdea7ffffffff"),
                (x"ffffffffff4801eed3bef7a619cfdeef7bdf5000053fffffff"),
                (x"ffffffffff65ee0053bef7bdef7bdef529d05ef7653fffffff"),
                (x"ffffffffff0318c0529def833087deed280bdef74b3fffffff"),
                (x"ffffffffff0318c0529def833087deed280bdef74b3fffffff"),
                (x"fffffffffff8000a5294a53bdef694a52804def74b3fffffff"),
                (x"fffffffffffffffa529def7deef7deef7b46252907ffffffff"),
                (x"fffffffffffffffa529defbdeef7beed294a0000ffffffffff"),
                (x"fffffffffffffffff39ce75ceef79ce738007fffffffffffff"),
                (x"fffffffffffffffff39ce75ceef79ce738007fffffffffffff"),
                (x"fffffffffffffffffc1deb9ae73bbce001ffffffffffffffff"),
                (x"fffffffffffffffffffce3bbdef41ce7ffffffffffffffffff"),
                (x"fffffffffffffffffffff80000001fffffffffffffffffffff"),

                -- 5_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffe94ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffe94a77ae739ad6b5ad73bbda7ffffffff"),
                (x"fffffffffffffffa77ae735ad6b5ad6b5ad6b5ceed3fffffff"),
                (x"fffffffffffffffa77ae735ad6b5ad6b5ad6b5ceed3fffffff"),
                (x"fffffffffffd29deb9ad6b5ad6b5ad6b5ad6b5ad753fffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b5ad777bda53fffffff"),
                (x"fffffffff4eb9ce6b9ad6b5ad6b5ae777bdefbbdeb3fffffff"),
                (x"fffffffff4eb9ce6b9ad6b5ad6b5ae777bdefbbdeb3fffffff"),
                (x"fffffffff4739ce735cd6b5ae73bbded29def5291f7fffffff"),
                (x"ffffffd29d739ce739ae739ddef69df77bdedef767ffffffff"),
                (x"ffffffd29d739ce739ce777b4ef7ddef7b7bdd2907ffffffff"),
                (x"ffffffd29deb9ce73bb4a53bdef7b7bdef7bdd8c67ffffffff"),
                (x"ffffff8014a77bda53bded3bdbdd2c63197bdd8cffffffffff"),
                (x"ffffff8014a77bda53bded3bdbdd2c63197bdd8cffffffffff"),
                (x"ffffffffe0f5294a53bde8c77bdd2500017bdc00ffffffffff"),
                (x"ffffffffff077bded28948d37bdd2400017bdc00ffffffffff"),
                (x"ffffffffffa319da5297b8d37bdee4ef7b7bdc00ffffffffff"),
                (x"ffffffffffa77b4ef694a3137bdee4f7bd7bdc00ffffffffff"),
                (x"ffffffffffa77b4ef694a3137bdee4f7bd7bdc00ffffffffff"),
                (x"fffffffffffd294eb3b4a5137bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffffffffa7694a5189bdef7bdef7ba400ffffffffff"),
                (x"ffffffffffffffffd294a528c4a6f7bdef7483ffffffffffff"),
                (x"ffffffffffffffffffbdef69d6318c6318007fffffffffffff"),
                (x"ffffffffffffffffffbdef69d6318c6318007fffffffffffff"),
                (x"fffffffffffffffff7bef7bb4a50000001ffffffffffffffff"),
                (x"ffffffffffffffff83def7bdda53a0e801dfffffffffffffff"),
                (x"ffffffffffffffff83bded3a0ef7a0a001dfffffffffffffff"),
                (x"fffffffffffffff07414a3194a51374801dfffffffffffffff"),
                (x"fffffffffffffff07414a3194a51374801dfffffffffffffff"),
                (x"fffffffffffffff0500c65ef4f7937b8000fffffffffffffff"),
                (x"fffffffffffffffed2894dee9f7a89b801dfffffffffffffff"),
                (x"fffffffffffffe0a7680026f7f7bd4077bdfffffffffffffff"),
                (x"fffffffffffffe0a53bde8000a501ca529dfffffffffffffff"),
                (x"fffffffffffffe0a53bde8000a501ca529dfffffffffffffff"),
                (x"fffffffffffffff07694a53bd0039def7bffffffffffffffff"),
                (x"fffffffffffffff073bdeb9dd0039de8000fffffffffffffff"),
                (x"ffffffffffffffff8000000000001fffffffffffffffffffff"),

                -- 5_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffff4eb9cd6b5ad6b5ad6b9dded294ffffffffff"),
                (x"ffffffffffa77ae6b5ad6b5ad6b5ad739ce777bded3fffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ae777ae73bbdef69ffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ae777ae73bbdef69ffffff"),
                (x"ffffffd29d739ce777bdefbdef7bdeed294a77bdef7b4a7fff"),
                (x"ffffffd29d739d4a77b4a77bdef7bded294a5294ef7b4a7fff"),
                (x"ffffffd294ef7bda77bdef58318d8cef7bded294ef7b4a7fff"),
                (x"ffffffd294ef7bda77bdef58318d8cef7bded294ef7b4a7fff"),
                (x"ffffff8014ed29deb19dea58318c6c4f7acef7bda768007fff"),
                (x"ffffffffe0ef7bdea6f7bdee918d37bdef7677bdef41ffffff"),
                (x"fffffffff403183edef7bdef7bdef7bdef7bf463e829ffffff"),
                (x"fffffffff460c6ceb2f7bdef7bdef7bdef76758c1f69ffffff"),
                (x"ffffffffffeb19d4a6f7bdef7bdef7bdef74a694677fffffff"),
                (x"ffffffffffeb19d4a6f7bdef7bdef7bdef74a694677fffffff"),
                (x"ffffffffffa319d4dd8c632f7bdef76318c4a694653fffffff"),
                (x"ffffffffff0529d4dca0002f7bdef700005ba694a03fffffff"),
                (x"ffffffffff05ef44dc80002f7bdef700004ba694b83fffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"ffffffffffffffd026f7bdef7bdef7bdef7483ffffffffffff"),
                (x"ffffffffffff7b4eb137bdef7bdef7bdee967694ef7fffffff"),
                (x"ffffffffffed29eed28c62537bdee94b19da77deed3bffffff"),
                (x"ffffffffffed29eed28c62537bdee94b19da77deed3bffffff"),
                (x"ffffffffe0a77bded3bded0e739ce7a77b4a7bdef77bffffff"),
                (x"ffffffffec6529da53bef7a80a5014f7bd4e8294e829deffff"),
                (x"fffffffbc94b180a53def7badef5bdf7bd40018cba41deffff"),
                (x"ffffffd29ef7bc0ed3def7a8def5b4f7bc065294a259ffffff"),
                (x"ffffffd29ef7bc0ed3def7a8def5b4f7bc065294a259ffffff"),
                (x"ffffffb194a52800769def81400280ef7acba694a03fffffff"),
                (x"ffffffb189bb180ed3b4a529def7bdef7acbdd29a03fffffff"),
                (x"ffffff80094801fed3def781d73ba0a52804dd2907ffffffff"),
                (x"ffffffffe00001f07694a501de73a0ef7bc00000ffffffffff"),
                (x"ffffffffe00001f07694a501de73a0ef7bc00000ffffffffff"),
                (x"ffffffffffffffff83bdeb9aeef41def39ffffffffffffffff"),
                (x"ffffffffffffffffff9deb9aeef41de801ffffffffffffffff"),
                (x"ffffffffffffffffffe00000000000ffffffffffffffffffff"),

                -- 5_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffdef7bdef7bda529fffffffffffffffffffff"),
                (x"ffffffffffa77ae735ad6b5ae73bbda529ffffffffffffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad777bda77ffffffffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad777bda77ffffffffffff"),
                (x"fffffffff4735ad6b5ad6b5ad6b5ad6b5aeef694ffffffffff"),
                (x"fffffffff4a77bd6b5ad6b5ad6b5ad6b5ad73bbda7ffffffff"),
                (x"ffffffffecef7beef7ae739ad6b5ad6b5ae6b9ceed3fffffff"),
                (x"ffffffffecef7beef7ae739ad6b5ad6b5ae6b9ceed3fffffff"),
                (x"fffffffffd1a53def69def7ae739ad6b9cd739ce753fffffff"),
                (x"ffffffffff65ef7ef7bef769def5ce735ae739ce7769ffffff"),
                (x"ffffffffff02537bdefdef7dda53bd739ce739ce7769ffffff"),
                (x"ffffffffff63197bdef7bdfbdef7b4a77ae739ceef69ffffff"),
                (x"fffffffffffb197bdd8c63137ef7b4ef7b4a77bda501ffffff"),
                (x"fffffffffffb197bdd8c63137ef7b4ef7b4a77bda501ffffff"),
                (x"fffffffffff8017bdc0001537bdc63ef7b4a5294f03fffffff"),
                (x"fffffffffff8017bdc0001137bdd234d29def7bd07ffffffff"),
                (x"fffffffffff8017bdfbde92f7bdd23bd294a758ca7ffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd2ca529ded3bda7ffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd2ca529ded3bda7ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a77aced294ffffffffff"),
                (x"fffffffffff8009bdef7bdef74a594a529da7fffffffffffff"),
                (x"fffffffffffffe04def7bdee963294a5294fffffffffffffff"),
                (x"fffffffffffffff0018c6318cef69def7bffffffffffffffff"),
                (x"fffffffffffffff0018c6318cef69def7bffffffffffffffff"),
                (x"fffffffffffffffffc0000014a53bef77bdfffffffffffffff"),
                (x"fffffffffffffffff41de83b4ef7def7bc0fffffffffffffff"),
                (x"fffffffffffffffff414a03bd003b4ef7a0fffffffffffffff"),
                (x"fffffffffffffffff4094dd34a518ca001d07fffffffffffff"),
                (x"fffffffffffffffff4094dd34a518ca001d07fffffffffffff"),
                (x"ffffffffffffffff8017bdd3ea52f76001407fffffffffffff"),
                (x"fffffffffffffffff417ba69e4a6f74d294effffffffffffff"),
                (x"fffffffffffffffff7a0053debdee90529da03ffffffffffff"),
                (x"fffffffffffffffff694a701400000ef7b4a03ffffffffffff"),
                (x"fffffffffffffffff694a701400000ef7b4a03ffffffffffff"),
                (x"fffffffffffffffffc1def780ef7b4a529d07fffffffffffff"),
                (x"ffffffffffffffff801def780ef5ceef7bc07fffffffffffff"),
                (x"fffffffffffffffffffffffe00000000000fffffffffffffff"),

                -- 5_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffff4ef5ce739ce739ce739ceef694ffffffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b9cd739ceed3fffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b9cd739ceed3fffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad6b5ae6b9ce7769ffffff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad739ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad735ce739d4a7fff"),
                (x"ffffffd28e6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4a7fff"),
                (x"ffffffd29d735ad6b5ad6b5ad6b5ad6b5ad735ce6bbb4a7fff"),
                (x"ffffffd29deb9ce6b5ad6b5ad6b5ad6b5ad6b9ad777b4a7fff"),
                (x"ffffffd294ef7bd739cd6b5ad6b5ad6b5ad73bbdef694a7fff"),
                (x"ffffffd294ef7bd739cd6b5ad6b5ad6b5ad73bbdef694a7fff"),
                (x"fffffffff4ef7bdef7ae739ce739ce739ddef7bdef69ffffff"),
                (x"ffffffffffa529def7bdef7bdef7bdef7bdef7bded3bffffff"),
                (x"ffffffffffef7b4a53bdef7bdef7bdef7bda5294ef7fffffff"),
                (x"ffffffffffff7bda5294a53bdef7bda5294a53bdefffffffff"),
                (x"ffffffffffff7bda5294a53bdef7bda5294a53bdefffffffff"),
                (x"fffffffffffffe0a77b4a77bdef7bded29def400ffffffffff"),
                (x"fffffffffffffff053ac653bdef7bdef7aca03ffffffffffff"),
                (x"ffffffffffffff4a529ded3b4ef69da5294a7694a7ffffffff"),
                (x"fffffffffffd294f7bb4a0294a5294a5294efbdea53fffffff"),
                (x"fffffffffffd294f7bb4a0294a5294a5294efbdea53fffffff"),
                (x"fffffffffffd29ef7bb4a5014a5294efbdda7bdef03fffffff"),
                (x"ffffffffffa0000a7bbdef7de9cc33f7bdda77de027fffffff"),
                (x"ffffffffffa3197b83b4a7bdef7bdef7bdda0000bb3fffffff"),
                (x"ffffffffff62537bdc14a77de08661f77b4a018c603fffffff"),
                (x"ffffffffff62537bdc14a77de08661f77b4a018c603fffffff"),
                (x"ffffffffff62537ba414a5294ef7bda5294a500007ffffffff"),
                (x"fffffffffff80094b29def7deef7deef7b4a53ffffffffffff"),
                (x"fffffffffffffe005294a77ddef7def77b4a53ffffffffffff"),
                (x"ffffffffffffffff801ce739cef5ceef39ce7fffffffffffff"),
                (x"ffffffffffffffff801ce739cef5ceef39ce7fffffffffffff"),
                (x"ffffffffffffffffffe00739d739cd777a0fffffffffffffff"),
                (x"ffffffffffffffffffffff380ef7bd7739ffffffffffffffff"),
                (x"fffffffffffffffffffffffe000000e7ffffffffffffffffff"),

                -- 5_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffe94ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffe94a77ae739ad6b5ad73bbda7ffffffff"),
                (x"fffffffffffffffa77ae735ad6b5ad6b5ad6b5ceed3fffffff"),
                (x"fffffffffffffffa77ae735ad6b5ad6b5ad6b5ceed3fffffff"),
                (x"fffffffffffd29deb9ad6b5ad6b5ad6b5ad6b5ad753fffffff"),
                (x"ffffffffffa77ae735ad6b5ad6b5ad6b5ad777bda53fffffff"),
                (x"fffffffff4eb9ce6b9ad6b5ad6b5ae777bdefbbdeb3fffffff"),
                (x"fffffffff4eb9ce6b9ad6b5ad6b5ae777bdefbbdeb3fffffff"),
                (x"fffffffff4739ce735cd6b5ae73bbded29def5291bffffffff"),
                (x"ffffffd29d739ce739ae739ddef69df77bdedef767ffffffff"),
                (x"ffffffd29d739ce739ce777b4ef7deef7b7bdd2907ffffffff"),
                (x"ffffffd29deb9ce73bb4a53bdef7bdbdef7bdd8c67ffffffff"),
                (x"ffffff8014a77bda53bded3bdbdd2c63197bdd8cffffffffff"),
                (x"ffffff8014a77bda53bded3bdbdd2c63197bdd8cffffffffff"),
                (x"ffffffffe0f5294a53bdef477bdd2500017bdc00ffffffffff"),
                (x"ffffffffff077bdef68948d37bdd2400017bdc00ffffffffff"),
                (x"ffffffffffa319da5297b8d37bdee4ef7b7bdc00ffffffffff"),
                (x"ffffffffffa77b4ef694a3137bdee4f7bd7bdc00ffffffffff"),
                (x"ffffffffffa77b4ef694a3137bdee4f7bd7bdc00ffffffffff"),
                (x"fffffffffffd294eb3b4a5137bdef7bdef7bdc00ffffffffff"),
                (x"fffffffffffffffa7694a5189bdef7bdef7ba400ffffffffff"),
                (x"ffffffffffffffffd294a768c4a6f7bdef7483ffffffffffff"),
                (x"fffffffffffffffef7dded3b439ce739ce007fffffffffffff"),
                (x"fffffffffffffffef7dded3b439ce739ce007fffffffffffff"),
                (x"ffffffffffffffdefbdef77deef41d077a0fffffffffffffff"),
                (x"ffffffffffffff4a77bef53def781d077a0a7fffffffffffff"),
                (x"fffffffffffffe003194a77bef7a8da35a067fffffffffffff"),
                (x"fffffffffffffe04a5200769df7a8da77b44b3ffffffffffff"),
                (x"fffffffffffffe04a5200769df7a8da77b44b3ffffffffffff"),
                (x"fffffffffffffe04dd3ef7a9def69da5280483ffffffffffff"),
                (x"fffffffffffffe06269ef5129a5294ef7a007fffffffffffff"),
                (x"fffffffffffffff0329ef52f7003bea77bdfffffffffffffff"),
                (x"fffffffffffffffef414a52f7003bda77bdfffffffffffffff"),
                (x"fffffffffffffffef414a52f7003bda77bdfffffffffffffff"),
                (x"fffffffffffffff003bded294a5294ef380fffffffffffffff"),
                (x"fffffffffffffffff39ce739def5c00739ffffffffffffffff"),
                (x"ffffffffffffffff839ce7c000001ce0000fffffffffffffff"),

                -- 5_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffd294a77bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffff4eb9cd6b5ad6b5ad6b9dded294ffffffffff"),
                (x"ffffffffffa77ae6b5ad6b5ad6b5ad739ce777bded3fffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ae777ae73bbdef69ffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ae777ae73bbdef69ffffff"),
                (x"ffffffd29d739ce777bdefbdef7bdeed294a77bdef7b4a7fff"),
                (x"ffffffd29d739d4a77b4a77bdef7bded294a5294ef7b4a7fff"),
                (x"ffffffd294ef7bda77bdef58318d8cef7bded294ef7b4a7fff"),
                (x"ffffffd294ef7bda77bdef58318d8cef7bded294ef7b4a7fff"),
                (x"ffffff8014ed29deb19dea58318c6c4f7acef7bda768007fff"),
                (x"ffffffffe0ef7bdea6f7bdee918d37bdef7677bdef41ffffff"),
                (x"fffffffff403183edef7bdef7bdef7bdef7bf463e829ffffff"),
                (x"fffffffff460c6ceb2f7bdef7bdef7bdef76758c1f69ffffff"),
                (x"ffffffffffeb19d4a6f7bdef7bdef7bdef74a694677fffffff"),
                (x"ffffffffffeb19d4a6f7bdef7bdef7bdef74a694677fffffff"),
                (x"ffffffffffa319d4dd8c632f7bdef76318c4a694653fffffff"),
                (x"ffffffffff0529d4dca0002f7bdef700005ba694a03fffffff"),
                (x"ffffffffff05ef44dc80002f7bdef700004ba694b83fffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffff80004dc9def6f7bdef7ef7a4ba40007ffffffff"),
                (x"fffffffffffffe065c9ef7af7bdef7f7bc4bb000ffffffffff"),
                (x"fffffffffffffff026f7bdef7bdef7bdef7483bdffffffffff"),
                (x"ffffffffffef7b4eb137bdef7bdef7bdee967694efffffffff"),
                (x"fffffffffda77beed3ac62537bdee94b194a77dea77fffffff"),
                (x"fffffffffda77beed3ac62537bdee94b194a77dea77fffffff"),
                (x"fffffffffdefbdef529ded0e739ce7a77bda77bded01ffffff"),
                (x"fffffff7b4077b40769ef7a80a5014f7bdda53bda319ffffff"),
                (x"fffffff7a04deec0029ef7badef5bdf7bdea50006252c67fff"),
                (x"ffffffffec4d294a301ef7a8def5b4f7bdea7400f7bcc67fff"),
                (x"ffffffffec4d294a301ef7a8def5b4f7bdea7400f7bcc67fff"),
                (x"ffffffffff052944dd9def41400280f77b4e8000a529ffffff"),
                (x"ffffffffff05289bdd9def7bdef7b4a529da740065d3ffffff"),
                (x"fffffffffff8009ba414a501d73ba0f7bdea77ff0253ffffff"),
                (x"fffffffffffffe00039def41de73a0a5294e83ff0001ffffff"),
                (x"fffffffffffffe00039def41de73a0a5294e83ff0001ffffff"),
                (x"fffffffffffffffffffce77a0ef5cd777bd07fffffffffffff"),
                (x"ffffffffffffffffffe0077a0ef5cd777bcfffffffffffffff"),
                (x"ffffffffffffffffffffffc00e70000001ffffffffffffffff"),

                -- 5_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffdef7bdef7bda529fffffffffffffffffffff"),
                (x"ffffffffffa77ae735ad6b5ae73bbda529ffffffffffffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad777bda7fffffffffffff"),
                (x"fffffffff4eb9cd6b5ad6b5ad6b5ad777bda7fffffffffffff"),
                (x"fffffffff4735ad6b5ad6b5ad6b5ad6b5aeef694ffffffffff"),
                (x"fffffffff4a77bd735ad6b5ad6b5ad6b5ad73bbda7ffffffff"),
                (x"ffffffffecef7beef7ae739ad6b5ad6b5ae6b9ceed3fffffff"),
                (x"ffffffffecef7beef7ae739ad6b5ad6b5ae6b9ceed3fffffff"),
                (x"fffffffffd1a53def69def7ae739ad6b9cd739ce753fffffff"),
                (x"ffffffffff65ef7ef7bef769def5ce735ae739ce7769ffffff"),
                (x"ffffffffff02537bdfbdef7dda53bd739ce739ce7769ffffff"),
                (x"ffffffffff63197bdef7bdfbdef7b4a77ae739ceef69ffffff"),
                (x"fffffffffffb197bdd8c63137ef7b4ef7b4a77bda501ffffff"),
                (x"fffffffffffb197bdd8c63137ef7b4ef7b4a77bda501ffffff"),
                (x"fffffffffff8017bdc0001537bdc63ef7b4a5294f03fffffff"),
                (x"fffffffffff8017bdc0001137bdd234d294ef7bd07ffffffff"),
                (x"fffffffffff8017bdfbde92f7bdd23bd294a758ca7ffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd2ca529ded3bda7ffffffff"),
                (x"fffffffffff8017bdfdef12f7bdd2ca529ded3bda7ffffffff"),
                (x"fffffffffff8017bdef7bdef7bdd34a77aced294ffffffffff"),
                (x"fffffffffff8009bdef7bdef74a594a529da7fffffffffffff"),
                (x"fffffffffffffe04def7bdee96329da5294fffffffffffffff"),
                (x"fffffffffffffff0018c6318ca53b4efbddeffffffffffffff"),
                (x"fffffffffffffff0018c6318ca53b4efbddeffffffffffffff"),
                (x"ffffffffffffffff83a00741df7bddf7bdeef7ffffffffffff"),
                (x"fffffffffffffffa03a00741ef7bd4f77bda53ffffffffffff"),
                (x"fffffffffffffff601b4a369ef7bbda318c003ffffffffffff"),
                (x"fffffffffffffec4d3b4a369eef69d02529483ffffffffffff"),
                (x"fffffffffffffec4d3b4a369eef69d02529483ffffffffffff"),
                (x"fffffffffffffe048294a769def69ef2537483ffffffffffff"),
                (x"fffffffffffffff003bded2944a534f5289603ffffffffffff"),
                (x"fffffffffffffffff7b4a7ba0bdef4f528c07fffffffffffff"),
                (x"fffffffffffffffff7b4a77a0bdef4a001deffffffffffffff"),
                (x"fffffffffffffffff7b4a77a0bdef4a001deffffffffffffff"),
                (x"ffffffffffffffff839ded294a5294ef7a007fffffffffffff"),
                (x"ffffffffffffffffff8e739ddef79ce739cfffffffffffffff"),
                (x"ffffffffffffffff8000000000001fe7380fffffffffffffff"),

                -- 6_character_0_0
                (x"fffffffffffffffffd8c677bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffffd8c677bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffa53bef787eef7def77bd633ffffffffffff"),
                (x"fffffffffffd29df7bddef863f787ef77b4ef7bda7ffffffff"),
                (x"ffffffffffa77be18fdef786318c7ef529da77deed3fffffff"),
                (x"ffffffffffa529df0c7ef77c318c7eed294efbbda53fffffff"),
                (x"ffffffffffa529df0c7ef77c318c7eed294efbbda53fffffff"),
                (x"ffffffffe0ef7b4ef87ef77c3f787eed29df7694ef69ffffff"),
                (x"ffffffffe0a7bdda77bef7bbeef47da529ded3bdf501ffffff"),
                (x"ffffffffe0a77beed29defbbeef7dda77bda03deed01ffffff"),
                (x"ffffffffe0a77beed29defbbeef7dda77bda03deed01ffffff"),
                (x"ffffffffe0ed29df7694a77bda53b4a77b4053bda501ffffff"),
                (x"ffffffffe0a77b4a7694a529da53b4a5294a5000a001ffffff"),
                (x"ffffffffff077bded294a5294a5294a5294a0294a03fffffff"),
                (x"ffffffffff0529def694a7694a5294a529405294003fffffff"),
                (x"ffffffffff0529def7b4a7694a5294a5294a5000003fffffff"),
                (x"ffffffffff0529def7b4a7694a5294a5294a5000003fffffff"),
                (x"ffffffffff0529df77bdef7b4a53b4a5294a0294003fffffff"),
                (x"ffffffffffa77bdf53bdefbb4ef7b4a77b4a5294a03fffffff"),
                (x"ffffffffffa77bdf53bdefbbdef7dda77b4a5000a03fffffff"),
                (x"ffffffffffefbddefa9defbb4ef7dda529da5000a03fffffff"),
                (x"ffffffffffefbddefa9defbb4ef7dda529da5000a03fffffff"),
                (x"ffffffffffefbd4ef81defbd4f7bdda529da5000a03fffffff"),
                (x"ffffffffffa77a0ef81defbd4f7bdd0529da5000a03fffffff"),
                (x"ffffffffff05280a7414a77c0ef7d40529d05000027fffffff"),
                (x"ffffffffe60528005014a77a0a53b405294050004a4dffffff"),
                (x"ffffffffe60528005014a77a0a53b405294050004a4dffffff"),
                (x"fffffffffe480090020005280a528005280001294a7dffffff"),
                (x"ffffffffec4b18cf01e528005000052800f0798c6259ffffff"),
                (x"ffffffffe04dee9077cf7c205294b083dfee8129ba41ffffff"),
                (x"ffffffffff00000677bdef8c6318c6f77bdeb000003fffffff"),
                (x"ffffffffff00000677bdef8c6318c6f77bdeb000003fffffff"),
                (x"fffffffffffffff074e73bde7ef4ef79ce7e83ffffffffffff"),
                (x"fffffffffffffffff4e73bde7ef4ef79ce7effffffffffffff"),
                (x"fffffffffffffffff7a739cfdef7a739cfdeffffffffffffff"),
                (x"ffffffffffffffff83bdef7bd003bdef7bd07fffffffffffff"),
                (x"ffffffffffffffff83bdef7bd003bdef7bd07fffffffffffff"),
                (x"ffffffffffffffff83bde9fbd003bd3f7bd07fffffffffffff"),
                (x"fffffffffffffffffc0739ce0ffc0739ce0fffffffffffffff"),
                (x"fffffffffffffffffc1defba0ffc1df77a0fffffffffffffff"),

                -- 6_character_0_1
                (x"fffffffffffffffffe94a77bdef694ef7ac633ffffffffffff"),
                (x"fffffffffffffffffe94a77bdef694ef7ac633ffffffffffff"),
                (x"fffffffffffffffa77bdef7def7bdea0c7eef694a7ffffffff"),
                (x"ffffffffffffff4ef694a77bdef463f77a3f0fbded3fffffff"),
                (x"fffffffffffd29da77bef7bdeef7be1fbde18fbdf77fffffff"),
                (x"ffffffffff05294ef7dded294a529df0c7e1fbbd1f7fffffff"),
                (x"ffffffffff05294ef7dded294a529df0c7e1fbbd1f7fffffff"),
                (x"ffffffffff0529def694a5289bdee9ed29df7694f53fffffff"),
                (x"ffffffffe0a5294a53bdef537bdef7bdef4ef529efffffffff"),
                (x"ffffffffe0a529def7b4a5137bdef7bdef7bdef767ffffffff"),
                (x"ffffffffe0a529def7b4a5137bdef7bdef7bdef767ffffffff"),
                (x"ffffffffe0a5294a0294a5137bdd9d4def7bdd2907ffffffff"),
                (x"ffffffffe0a00000529def5374a534ef7a9bdd8ca7ffffffff"),
                (x"ffffffffe0a77b4a53bded3b7bdd2ca529dbde94ffffffffff"),
                (x"ffffffffe0a77b4ed3b4a7697bdee500009bdc00ffffffffff"),
                (x"ffffffffe0a77b4ed294a7a97bdee400017bdc00ffffffffff"),
                (x"ffffffffe0a77b4ed294a7a97bdee400017bdc00ffffffffff"),
                (x"fffffffff4ed29da501defa97bdee4e7397bdc00ffffffffff"),
                (x"fffffffff4e801d0501defa97bdee4739d7bdc00ffffffffff"),
                (x"fffffffff4a001d0501defa97bdef7bdef7bdc00ffffffffff"),
                (x"fffffffff4a001400014a7a89bdef7bdef7ba400ffffffffff"),
                (x"fffffffff4a001400014a7a89bdef7bdef7ba400ffffffffff"),
                (x"ffffffffe0a000000294a758c4a6f7bdef7483ffffffffffff"),
                (x"ffffffffe0a0000003c00519e6318c6318007fffffffffffff"),
                (x"ffffffffe0a000007929482067bcc66001efffffffffffffff"),
                (x"ffffffffe000000f26e9498cff78a587bcff7fffffffffffff"),
                (x"ffffffffe000000f26e9498cff78a587bcff7fffffffffffff"),
                (x"ffffffffff00000f5ee94a526f7bc58421ef7fffffffffffff"),
                (x"ffffffffffffffff5efef798c0001e84210f7fffffffffffff"),
                (x"fffffffffffffff05ef7bdd37bdd20294b0f7fffffffffffff"),
                (x"fffffffffffffff032f7bdef7bdee0814aff7fffffffffffff"),
                (x"fffffffffffffff032f7bdef7bdee0814aff7fffffffffffff"),
                (x"ffffffffffffffff8137bdd37bdd20318defffffffffffffff"),
                (x"fffffffffffffffffc000318c000c6318dffffffffffffffff"),
                (x"fffffffffffffffffc1def7bdef4e7ed29ffffffffffffffff"),
                (x"ffffffffffffffffffe0077bd39de7a7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0077bd39de7a7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0077a77bcfdffffffffffffffffffff"),
                (x"fffffffffffffffffffff83af7bde0ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83be297c0ffffffffffffffffffff"),

                -- 6_character_0_2
                (x"fffffffffffffffffe94a77bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffffe94a77bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffa53bdef87eef7def77bda53ffffffffffff"),
                (x"fffffffffffd29df769ef7463f787eef7b4ef7bda7ffffffff"),
                (x"ffffffffffa77be1fbb4a7ba318c7eed29da77deed3fffffff"),
                (x"ffffffffffa529df0fddefbbe18fdda5294efbbda53fffffff"),
                (x"ffffffffffa529df0fddefbbe18fdda5294efbbda53fffffff"),
                (x"ffffffffe0ef7b4e8fb4a53bdf7bbda529df7694ef41ffffff"),
                (x"ffffffffe0a7bdda7537ba69def7b44dee9a53bdf501ffffff"),
                (x"ffffffffe0a77bea5ef7bdee9ef537bdef7bd3deed01ffffff"),
                (x"ffffffffe0a77bea5ef7bdee9ef537bdef7bd3deed01ffffff"),
                (x"ffffffffe0a001da5ef7bdef7bdef7bdef7bd3bda501ffffff"),
                (x"ffffffffe0a77a0a33a94def7bdef7ba53d65294ed01ffffff"),
                (x"ffffffffffa77b44a69def537bdee9ef7b44a400ed3fffffff"),
                (x"ffffffffff077beea594a53b7bdefda528c4d3bda03fffffff"),
                (x"ffffffffff077bea5ca000137bdee900005bd3dea03fffffff"),
                (x"ffffffffff077bea5ca000137bdee900005bd3dea03fffffff"),
                (x"ffffffffff0529ea5c80002f7bdef700004bd3dea03fffffff"),
                (x"ffffffffffa529d05c9ce72f7bdef7e7384bd3dea53fffffff"),
                (x"ffffffffffa001d05c8e73af7bdef7739c4b83bd053fffffff"),
                (x"ffffffffffe801d026f7bdef7bdef7bdef7483bd077fffffff"),
                (x"ffffffffffe801d026f7bdef7bdef7bdef7483bd077fffffff"),
                (x"ffffffffff3001403137bdef7bdef7bdee96029401bfffffff"),
                (x"ffffffffe64a53403ccc62537bdee94b186782944a4dffffff"),
                (x"ffffff98c94a52603de52998c6318c314af780c64a52637fff"),
                (x"fffff3253ef252933de5294be4a7c52c20f799294fbc949bff"),
                (x"fffff3253ef252933de5294be4a7c52c20f799294fbc949bff"),
                (x"fffff331894b189f0205294aff79e5294b0079296252c61bff"),
                (x"fffff62537ba52c00205294a5294a5294b00018c4dee94b3ff"),
                (x"fffff625374def7600c5294a5294a5294a6032f7ba6e94b3ff"),
                (x"ffffff80094def7677c63421084210818deeb2f7ba52007fff"),
                (x"ffffff80094def7677c63421084210818deeb2f7ba52007fff"),
                (x"ffffffffe04def7074fef7bc6318def7bc7e82f7ba41ffffff"),
                (x"ffffffffff00000ff4e73bdef7bdef79ce7efc00003fffffff"),
                (x"ffffffffffffffffd3a73bcfda53a779cfda7fffffffffffff"),
                (x"ffffffffffffffff83a739cfd003a739cfd07fffffffffffff"),
                (x"ffffffffffffffff83a739cfd003a739cfd07fffffffffffff"),
                (x"ffffffffffffffff83af7bcfd003a77bdfd07fffffffffffff"),
                (x"fffffffffffffffffc1def7a0ffc1def7a0fffffffffffffff"),
                (x"ffffffffffffffffffbdefba0ffc1df77bdfffffffffffffff"),

                -- 6_character_0_3
                (x"ffffffffffffff4a53bded29def7bda529ffffffffffffffff"),
                (x"ffffffffffffff4a53bded29def7bda529ffffffffffffffff"),
                (x"ffffffffffa529def874a7bdef7bddef7bda7fffffffffffff"),
                (x"fffffffff4ef7a3f0fbef0c7def7bda529ded3ffffffffffff"),
                (x"fffffffffdf77a31fbc31fbbdf7bdef77bda7694ffffffffff"),
                (x"fffffffffd1f7be1f87ef7694a5294efbdded29407ffffffff"),
                (x"fffffffffd1f7be1f87ef7694a5294efbdded29407ffffffff"),
                (x"fffffffff4f529df769dea6f74a694a529def69407ffffffff"),
                (x"ffffffffffea53ded2f7bdef7bdd3def7b4a5294a03fffffff"),
                (x"ffffffffff65ef7bdef7bdef7bdd34a77bdef694a03fffffff"),
                (x"ffffffffff65ef7bdef7bdef7bdd34a77bdef694a03fffffff"),
                (x"ffffffffff02537bdee94f597bdd34a5280a5294a03fffffff"),
                (x"ffffffffffa3197ba7bded129bdd3ded29400000a03fffffff"),
                (x"fffffffffffd297bf694a3137bdfb4ef7b4a53bda03fffffff"),
                (x"fffffffffff8017ba400016f7bde9da77b4ed3bda03fffffff"),
                (x"fffffffffff8017bdc00012f7bde9ea5294ed3bda03fffffff"),
                (x"fffffffffff8017bdc00012f7bde9ea5294ed3bda03fffffff"),
                (x"fffffffffff8017bdf9ce12f7bde9ee8014a7694ed3fffffff"),
                (x"fffffffffff8017bddce712f7bde9ee801407400ed3fffffff"),
                (x"fffffffffff8017bdef7bdef7bde9ee801407400a53fffffff"),
                (x"fffffffffff8009bdef7bdef74a69ea000005000a53fffffff"),
                (x"fffffffffff8009bdef7bdef74a69ea000005000a53fffffff"),
                (x"fffffffffffffe04def7bdee96319da528000000a03fffffff"),
                (x"fffffffffffffff0018c6318cf799407bc000000a03fffffff"),
                (x"fffffffffffffffff80c618cf319204a53e00000a03fffffff"),
                (x"ffffffffffffffff3fd0814be7bd264dee9f0000003fffffff"),
                (x"ffffffffffffffff3fd0814be7bd264dee9f0000003fffffff"),
                (x"ffffffffffffffff7a10817de319294def7f000007ffffffff"),
                (x"ffffffffffffffff3cb0878006319ebdef7f7fffffffffffff"),
                (x"ffffffffffffffff40a528137bdd37bdef707fffffffffffff"),
                (x"ffffffffffffffff3cb0802f7bdef7bdeec07fffffffffffff"),
                (x"ffffffffffffffff3cb0802f7bdef7bdeec07fffffffffffff"),
                (x"ffffffffffffffff98c630137bdd37ba520fffffffffffffff"),
                (x"fffffffffffffffffe86318006318c0001ffffffffffffffff"),
                (x"fffffffffffffffffe9de9cfdef7bde801ffffffffffffffff"),
                (x"fffffffffffffffffff4a1de7ef7bd07ffffffffffffffffff"),
                (x"fffffffffffffffffff4a1de7ef7bd07ffffffffffffffffff"),
                (x"ffffffffffffffffffffff4ef39fbd07ffffffffffffffffff"),
                (x"fffffffffffffffffffff81ef7bfa0ffffffffffffffffffff"),
                (x"fffffffffffffffffffff83c5f7ba0ffffffffffffffffffff"),

                -- 6_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffa53bef787eef7def77bda53ffffffffffff"),
                (x"fffffffffffd29df7bddef863f787ef77b4ef7bda7ffffffff"),
                (x"ffffffffffa77be18fdef786318c7ef529da77deed3fffffff"),
                (x"ffffffffffa77be18fdef786318c7ef529da77deed3fffffff"),
                (x"ffffffffffa529df0c7ef77c318c7eed294efbbda53fffffff"),
                (x"ffffffffe0ef7b4ef87ef77c3f787eed29df7694ef69ffffff"),
                (x"ffffffffe0a7bdda77bef7bbeef47da529ded3bdf501ffffff"),
                (x"ffffffffe0a7bdda77bef7bbeef47da529ded3bdf501ffffff"),
                (x"ffffffffe0a77beed29defbbeef7dda77bda03deed01ffffff"),
                (x"ffffffffe0ed29df7694a77bda53b4a77b4053bda501ffffff"),
                (x"ffffffffe0a77b4a7694a529da53b4a5294a5000a001ffffff"),
                (x"ffffffffff077bded294a5294a5294a5294a0294a03fffffff"),
                (x"ffffffffff0529def7b4a7694a5294a529405294003fffffff"),
                (x"ffffffffff0529def7b4a7694a5294a529405294003fffffff"),
                (x"ffffffffff0529def7b4a7694a5294a5294a52940001ffffff"),
                (x"ffffffffff0529ef77d4a77b4a53b4a5294a5000a001ffffff"),
                (x"ffffffffff077beed3d4a77b4a53b4a5294a5294a001ffffff"),
                (x"ffffffffffa77bea77ddef7bda53bda5294a5294a501ffffff"),
                (x"ffffffffffa77bea77ddef7bda53bda5294a5294a501ffffff"),
                (x"ffffffffffa77bea77ddef7bda53bded294a52940501ffffff"),
                (x"fffffffffffd29d077d4a7bdda53beed294052940501ffffff"),
                (x"fffffffffff529d053b4a77dda53bee8014052940501ffffff"),
                (x"fffffffffff001400280053d4a529ee801405294003fffffff"),
                (x"fffffffffff001400280053d4a529ee801405294003fffffff"),
                (x"fffffffffff252080000053b40029da0014050004fbfffffff"),
                (x"ffffffffff67bdef1a05282940029404200781294fbfffffff"),
                (x"ffffffffff0318c019f081400294007bde64a529f33fffffff"),
                (x"fffffffffff8000078cf7be107bdfef7bc0f7bde4b3fffffff"),
                (x"fffffffffff8000078cf7be107bdfef7bc0f7bde4b3fffffff"),
                (x"ffffffffffffffffd0c6318c6318c6318d46252907ffffffff"),
                (x"ffffffffffffffffd3bde9defef7a73f7b4a0000ffffffffff"),
                (x"ffffffffffffffffd29def4e7ef694a528007fffffffffffff"),
                (x"fffffffffffffffffc14a77bd39c1de801ffffffffffffffff"),
                (x"fffffffffffffffffc14a77bd39c1de801ffffffffffffffff"),
                (x"ffffffffffffffffffe0050e7a500007ffffffffffffffffff"),
                (x"fffffffffffffffffffff83c3f781fffffffffffffffffffff"),
                (x"fffffffffffffffffffff83ddef41fffffffffffffffffffff"),

                -- 6_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffd8c677bdef694ef7b4a53ffffffffffff"),
                (x"fffffffffffffff677bdef7def7bdea0c7eef694a7ffffffff"),
                (x"ffffffffffffff4ef694a77bdef463f77a3f0fbded3fffffff"),
                (x"fffffffffffd29da77bef7bdeef7be1fbde18fbdf77fffffff"),
                (x"fffffffffffd29da77bef7bdeef7be1fbde18fbdf77fffffff"),
                (x"ffffffffff05294ef7dded294a529df0c7e1fbbd1f7fffffff"),
                (x"ffffffffff0529def694a5289bdee9ed29df7694f53fffffff"),
                (x"ffffffffe0a5294a53bdef537bdef7bdef4ef529efffffffff"),
                (x"ffffffffe0a5294a53bdef537bdef7bdef4ef529efffffffff"),
                (x"ffffffffe0a529def7b4a5137bdef7bdef7bdef767ffffffff"),
                (x"ffffffffe0a5294a0294a5137bdd9d4def7bdd2907ffffffff"),
                (x"ffffffffe0a77b40529def5374a534ef7a9bdd8ca7ffffffff"),
                (x"ffffffffe0ed29da53bded3b7bdd2ca529dbde94ffffffffff"),
                (x"ffffff8014ed29da03b4a7697bdee500009bdc00ffffffffff"),
                (x"ffffff8014ed29da03b4a7697bdee500009bdc00ffffffffff"),
                (x"ffffff801da77bda0294a7a97bdee400017bdc00ffffffffff"),
                (x"ffffff801da77b40001defa97bdee4e7397bdc00ffffffffff"),
                (x"ffffff801da77b40001defbb7bdee4739d7bdc00ffffffffff"),
                (x"fffff0529da77b400014a7bb7bdef7bdef7bdc00ffffffffff"),
                (x"fffff0529da77b400014a7bb7bdef7bdef7bdc00ffffffffff"),
                (x"fffff05294ed28000014a77ccbdef7bdef7ba400ffffffffff"),
                (x"fffff05280ed28000280053ac4a6f7bdef7483ffffffffffff"),
                (x"ffffffd280a0000003c94828c6318c6318007fffffffffffff"),
                (x"ffffff8000a0000002f7ba409f78c63001efffffffffffffff"),
                (x"ffffff8000a0000002f7ba409f78c63001efffffffffffffff"),
                (x"ffffffffe00001f07af7ba52931a1087bcf07fffffffffffff"),
                (x"ffffffffff0001f07937bdd29f79f087bc607fffffffffffff"),
                (x"fffffffffffffff018d7bdefef7800018cff7fffffffffffff"),
                (x"fffffffffffffff01bc94dee9632f7b800ff7fffffffffffff"),
                (x"fffffffffffffff01bc94dee9632f7b800ff7fffffffffffff"),
                (x"fffffffffffffff078c0026f74a6f7b8006f7fffffffffffff"),
                (x"fffffffffffffffe83def01374a537677a0fffffffffffffff"),
                (x"fffffffffffffffef4e73f40c63000077bffffffffffffffff"),
                (x"fffffffffffffff074ef79fbd003bdefffffffffffffffffff"),
                (x"fffffffffffffff074ef79fbd003bdefffffffffffffffffff"),
                (x"fffffffffffffff077a73f7bd003a73f7bffffffffffffffff"),
                (x"ffffffffffffffff80ef79fa00001df7bdffffffffffffffff"),
                (x"ffffffffffffffff83bef17c0fffffffffffffffffffffffff"),

                -- 6_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffa53bdef87eef7def77bda53ffffffffffff"),
                (x"fffffffffffd29df769ef7463f787eef7b4ef7bda7ffffffff"),
                (x"ffffffffffa77be1fbb4a7ba318c7eed29da77deed3fffffff"),
                (x"ffffffffffa77be1fbb4a7ba318c7eed29da77deed3fffffff"),
                (x"ffffffffffa529df0fddefbbe18fdda5294efbbda53fffffff"),
                (x"ffffffffe0ef7b4e8fb4a53bdf7bbda529df7694ef41ffffff"),
                (x"ffffffffe0a7bdda7537ba69def7b44dee9a53bdf501ffffff"),
                (x"ffffffffe0a7bdda7537ba69def7b44dee9a53bdf501ffffff"),
                (x"ffffffffe0a77bea5ef7bdee9ef537bdef7bd3deed01ffffff"),
                (x"ffffffffe0a001da5ef7bdef7bdef7bdef7bd3bda501ffffff"),
                (x"ffffffffe0a77a0a33a94def7bdef7ba53d65294ed01ffffff"),
                (x"ffffffffffa77b44a69def537bdee9ef7b44a400ed3fffffff"),
                (x"ffffffffff077beea594a53b7bdefda528c4d3bda03fffffff"),
                (x"ffffffffff077beea594a53b7bdefda528c4d3bda03fffffff"),
                (x"ffffffffff077bea5ca000137bdee900005bd3dea03fffffff"),
                (x"ffffffffff0529ea5c80002f7bdef700004bd3dea03fffffff"),
                (x"ffffffffffa529d05c9ce72f7bdef7e7384bd3dea53fffffff"),
                (x"ffffffffffa001d05c8e73af7bdef7739c4b83bd0769ffffff"),
                (x"ffffffffffa001d05c8e73af7bdef7739c4b83bd0769ffffff"),
                (x"ffffffffffa001d026f7bdef7bdef7bdef7483bd0769ffffff"),
                (x"ffffffffff3001403137bdef7bdef7bdee96029407ba007fff"),
                (x"ffffffffe64a53403c0c62537bdee94b180302944a7c007fff"),
                (x"fffffffbc94a529040c52998c6318c34206781294a53ef7fff"),
                (x"fffffffbc94a529040c52998c6318c34206781294a53ef7fff"),
                (x"fffffffbc94a52933cc5294be4a7c52c206341294a53ef7fff"),
                (x"ffffffb1894a52901a05294aff79e5294b0301294a7dffffff"),
                (x"ffffffb1894a52c01a05294a5294a5294a0032f7ba59ffffff"),
                (x"ffffffb197ba520f99e5294a5294a52bdecbdef74a59ffffff"),
                (x"ffffffb197ba520f99e5294a5294a52bdecbdef74a59ffffff"),
                (x"ffffffb189bb180ff7c6318c6318c637bccbdd296301ffffff"),
                (x"ffffff80094b19fff4e73bdef7bce73f7a04dd8c003fffffff"),
                (x"ffffffffe00001fff7a73bde7ef7bdef7bd00000ffffffffff"),
                (x"ffffffffffffffffffa739de739c1def7bdfffffffffffffff"),
                (x"ffffffffffffffffffa739de739c1def7bdfffffffffffffff"),
                (x"fffffffffffffffffffdebdef39c1def7bffffffffffffffff"),
                (x"ffffffffffffffffffe0077bdef40007ffffffffffffffffff"),
                (x"ffffffffffffffffffffff7beef7ffffffffffffffffffffff"),

                -- 6_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffff4a53bded29def7bda529ffffffffffffffff"),
                (x"ffffffffffa529def874a7bdef7bddef7bda7fffffffffffff"),
                (x"fffffffff4ef7a3f0fbef0c7def7bda529ded3ffffffffffff"),
                (x"fffffffffdf77a31fbc31fbbdf7bdef77bda7694ffffffffff"),
                (x"fffffffffdf77a31fbc31fbbdf7bdef77bda7694ffffffffff"),
                (x"fffffffffd1f7be1f87ef7694a5294efbdded29407ffffffff"),
                (x"fffffffff4f529df769dea6f74a694a529def69407ffffffff"),
                (x"ffffffffffea53ded2f7bdef7bdd3def7b4a5294a03fffffff"),
                (x"ffffffffffea53ded2f7bdef7bdd3def7b4a5294a03fffffff"),
                (x"ffffffffff65ef7bdef7bdef7bdd34a77bdef694a03fffffff"),
                (x"ffffffffff02537bdee94f597bdd34a5280a5294a03fffffff"),
                (x"ffffffffffa3197ba7bded129bdd3ded294053bda03fffffff"),
                (x"fffffffffffd297bf694a3137bdfb4ef7b4a7694e83fffffff"),
                (x"fffffffffff8017ba400016f7bde9da77a0a7694ed01ffffff"),
                (x"fffffffffff8017ba400016f7bde9da77a0a7694ed01ffffff"),
                (x"fffffffffff8017bdc00012f7bde9ea5280a77bda741ffffff"),
                (x"fffffffffff8017bdf9ce12f7bde9ee8000053bda741ffffff"),
                (x"fffffffffff8017bddce712f7bdfbee8000053bda741ffffff"),
                (x"fffffffffff8017bdef7bdef7bdfbea0000053bda768007fff"),
                (x"fffffffffff8017bdef7bdef7bdfbea0000053bda768007fff"),
                (x"fffffffffff8009bdef7bdef7633dda000000294ed28007fff"),
                (x"fffffffffffffe04def7bdee9633b40528000294e828007fff"),
                (x"fffffffffffffff0018c6318c632804fbc000000a029ffffff"),
                (x"fffffffffffffffff806318de4a409ba52000000a001ffffff"),
                (x"fffffffffffffffff806318de4a409ba52000000a001ffffff"),
                (x"fffffffffffffff03e10843c64a537ba53e07c00003fffffff"),
                (x"fffffffffffffff01a10879fe4a537ba53e07c0007ffffffff"),
                (x"ffffffffffffffff3cc00001ef7af7b98c607fffffffffffff"),
                (x"ffffffffffffffff3c17bdeec4a6f74fbc607fffffffffffff"),
                (x"ffffffffffffffff3c17bdeec4a6f74fbc607fffffffffffff"),
                (x"ffffffffffffffff1817bdee9bdee9018de07fffffffffffff"),
                (x"ffffffffffffffff83ac65d29bdd20f7bc0effffffffffffff"),
                (x"ffffffffffffffffffa00000c6301d39cfdeffffffffffffff"),
                (x"fffffffffffffffffffdef7a0ef7a779cfd07fffffffffffff"),
                (x"fffffffffffffffffffdef7a0ef7a779cfd07fffffffffffff"),
                (x"ffffffffffffffffffa739fa0ef7bd3f7bd07fffffffffffff"),
                (x"ffffffffffffffffffdef7400003a779ce0fffffffffffffff"),
                (x"fffffffffffffffffffffffff003c5f77a0fffffffffffffff"),

                -- 6_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffa53bef787eef7def77bda53ffffffffffff"),
                (x"fffffffffffd29df7bddef863f787ef77b4ef7bda7ffffffff"),
                (x"ffffffffffa77be18fdef786318c7ef529da77deed3fffffff"),
                (x"ffffffffffa77be18fdef786318c7ef529da77deed3fffffff"),
                (x"ffffffffffa529df0c7ef77c318c7eed294efbbda53fffffff"),
                (x"ffffffffe0ef7b4ef87ef77c3f787eed29df7694ef69ffffff"),
                (x"ffffffffe0a7bdda77bef7bbeef47da529ded3bdf501ffffff"),
                (x"ffffffffe0a7bdda77bef7bbeef47da529ded3bdf501ffffff"),
                (x"ffffffffe0a77beed29defbbeef7dda77bda03deed01ffffff"),
                (x"ffffffffe0ed29df7694a77bda53b4a77b4053bda501ffffff"),
                (x"ffffffffe0a77b4a7694a529da53b4a5294a5000a001ffffff"),
                (x"ffffffffff077bded294a5294a5294a5294a0294a03fffffff"),
                (x"ffffffffff077bdef694a7694a5294a529405294003fffffff"),
                (x"ffffffffff077bdef694a7694a5294a529405294003fffffff"),
                (x"ffffffffffa77bdef694a77bda5294a5294a5000003fffffff"),
                (x"ffffffffffa77bdef69def7bda5294a5294a5294003fffffff"),
                (x"ffffffffffa77bdf769def7bda53b4a77b4a5294003fffffff"),
                (x"fffffffff4f77b4f769def7bda53b4a77b4a0294003fffffff"),
                (x"fffffffff4f77b4f769def7bda53b4a77b4a0294003fffffff"),
                (x"fffffffff4f529df769def41def7b4a77b4a029407ffffffff"),
                (x"fffffffffeed29eed3bef741df7bb4ef7b40529407ffffffff"),
                (x"fffffffffd0529ea53def501df7bb4ef7b40529407bfffffff"),
                (x"fffffffff400014053dded014f7a80ed294050004fbfffffff"),
                (x"fffffffff400014053dded014f7a80ed294050004fbfffffff"),
                (x"fffffffffff2520053dde8014ef680ed280a50004fbfffffff"),
                (x"fffffffffff2529483b4a0014a5000a0000003def33fffffff"),
                (x"ffffffffff67bc94a40003e00000a50000f3018c603fffffff"),
                (x"ffffffffff6253ef781ef7bcf7be107bde6f000007ffffffff"),
                (x"ffffffffff6253ef781ef7bcf7be107bde6f000007ffffffff"),
                (x"fffffffffff80094b29def7bdef4c6318c6a7fffffffffffff"),
                (x"fffffffffffffe00529de9cfdef5ef3f7bda7fffffffffffff"),
                (x"ffffffffffffffff8014a5294ef4e7ef7b4a7fffffffffffff"),
                (x"ffffffffffffffffffe0077a039fbded280fffffffffffffff"),
                (x"ffffffffffffffffffe0077a039fbded280fffffffffffffff"),
                (x"fffffffffffffffffffff8000a50e7a001ffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f787e07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0ef7be07ffffffffffffffffff"),

                -- 6_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bdef694ef7b4a53ffffffffffff"),
                (x"fffffffffffffffa77bdef7def7bdea0c7eef694a7ffffffff"),
                (x"ffffffffffffff4ef694a77bdef463f77a3f0fbded3fffffff"),
                (x"fffffffffffd29da77bef7bdeef7be1fbde18fbdf77fffffff"),
                (x"fffffffffffd29da77bef7bdeef7be1fbde18fbdf77fffffff"),
                (x"ffffffffff05294ef7dded294a529df0c7e1fbbd1f7fffffff"),
                (x"ffffffffff0529def694a5289bdee9ed29df7694f53fffffff"),
                (x"ffffffffe0a5294a53bdef537bdef7bdef4ef529efffffffff"),
                (x"ffffffffe0a5294a53bdef537bdef7bdef4ef529efffffffff"),
                (x"ffffffffe0a529def7b4a5137bdef7bdef7bdef767ffffffff"),
                (x"ffffffffe0a5294a5294a5137bdd9d4def7bdd2907ffffffff"),
                (x"ffffffffe00529da501def5374a534ef7a9bdd8ca7ffffffff"),
                (x"ffffffffe00529da53bded3b7bdd2ca529dbde94ffffffffff"),
                (x"ffffffffe0a529da53b4a7697bdee500009bdc00ffffffffff"),
                (x"ffffffffe0a529da53b4a7697bdee500009bdc00ffffffffff"),
                (x"ffffffffe0a77b4ed294a7a97bdee400017bdc00ffffffffff"),
                (x"fffffffff4a77b4ed01defa97bdee4e7397bdc00ffffffffff"),
                (x"fffffffff4a77b4a001defa97bdee4739d7bdc00ffffffffff"),
                (x"fffffffff4a77a0a001defa97bdef7bdef7bdc00ffffffffff"),
                (x"fffffffff4a77a0a001defa97bdef7bdef7bdc00ffffffffff"),
                (x"fffffffff4a77a000014a7a89bdef7bdef7ba400ffffffffff"),
                (x"ffffffffe0a77a000294a758c4a6f7bdef7483ffffffffffff"),
                (x"ffffffffe0a77a0001200519e6318c6318007fffffffffffff"),
                (x"ffffffffff05280026e9480cf840c64801efffffffffffffff"),
                (x"ffffffffff05280026e9480cf840c64801efffffffffffffff"),
                (x"ffffffffff05280f5ee94a5fe294b0f420ff7fffffffffffff"),
                (x"fffffffffff800035ee94a5ef8421087bcf67fffffffffffff"),
                (x"fffffffffffffe04def7ba7c68421083dfe4b3ffffffffffff"),
                (x"fffffffffffffe0f26f7ba4008421083dfe483ffffffffffff"),
                (x"fffffffffffffe0f26f7ba4008421083dfe483ffffffffffff"),
                (x"fffffffffffffff026f7bdee9f79ef7fbc007fffffffffffff"),
                (x"fffffffffffffff03137bdef7000c6318c0fffffffffffffff"),
                (x"ffffffffffffffff800c626e9001ef3f7bffffffffffffffff"),
                (x"ffffffffffffffff83bde8000ef4fdef7bffffffffffffffff"),
                (x"ffffffffffffffff83bde8000ef4fdef7bffffffffffffffff"),
                (x"fffffffffffffffff7bde8000ef4ef79cfffffffffffffffff"),
                (x"ffffffffffffffff801def400003a7ef7a0fffffffffffffff"),
                (x"fffffffffffffffffffffffff003be2fbc0fffffffffffffff"),

                -- 6_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bdef7bded294fffffffffffffff"),
                (x"fffffffffffffffa53bdef87eef7def77bda53ffffffffffff"),
                (x"fffffffffffd29df769ef7463f787eef7b4ef7bda7ffffffff"),
                (x"ffffffffffa77be1fbb4a7ba318c7eed29da77deed3fffffff"),
                (x"ffffffffffa77be1fbb4a7ba318c7eed29da77deed3fffffff"),
                (x"ffffffffffa529df0fddefbbe18fdda5294efbbda53fffffff"),
                (x"ffffffffe0ef7b4e8fb4a53bdf7bbda529df7694ef41ffffff"),
                (x"ffffffffe0a7bdda7537ba69def7b44dee9a53bdf501ffffff"),
                (x"ffffffffe0a7bdda7537ba69def7b44dee9a53bdf501ffffff"),
                (x"ffffffffe0a77bea5ef7bdee9ef537bdef7bd3deed01ffffff"),
                (x"ffffffffe0a001da5ef7bdef7bdef7bdef7bd3bda501ffffff"),
                (x"ffffffffe0a77a0a33a94def7bdef7ba53d65294ed01ffffff"),
                (x"ffffffffffa77b44a69def537bdee9ef7b44a400ed3fffffff"),
                (x"ffffffffff077beea594a53b7bdefda528c4d3bda03fffffff"),
                (x"ffffffffff077beea594a53b7bdefda528c4d3bda03fffffff"),
                (x"ffffffffff077bea5ca000137bdee900005bd3dea03fffffff"),
                (x"ffffffffff0529ea5c80002f7bdef700004bd3dea03fffffff"),
                (x"fffffffff4a529d05c9ce72f7bdef7e7384bd3dea53fffffff"),
                (x"fffffffff4e801d05c8e73af7bdef7739c4b83bd053fffffff"),
                (x"fffffffff4e801d05c8e73af7bdef7739c4b83bd053fffffff"),
                (x"fffffffff4e801d026f7bdef7bdef7bdef7483bd053fffffff"),
                (x"ffffffd29df001403137bdef7bdef7bdee96029401bfffffff"),
                (x"fffffffbde4a5340180c62537bdee94b180782944a4dffffff"),
                (x"fffffffbc94a52903cd08198c6318c314a6801294a53ef7fff"),
                (x"fffffffbc94a52903cd08198c6318c314a6801294a53ef7fff"),
                (x"fffffffbc94a529498d0814be4a7c52c206799294a53ef7fff"),
                (x"fffffffbc94a52901a05294aff79e5294b0301294b12c67fff"),
                (x"ffffffffec4def760005294a5294a5294b03018c6252c67fff"),
                (x"ffffffffec4a537bdd8f794a5294a5294af37c004deec67fff"),
                (x"ffffffffec4a537bdd8f794a5294a5294af37c004deec67fff"),
                (x"ffffffffe063189bdd9ef18c6318c67fbdeefc0065d2c67fff"),
                (x"ffffffffff0000cba41de9ce77bdef79ce7effff6252007fff"),
                (x"fffffffffffffe0003bdef7bdef4ef79cfdeffff0001ffffff"),
                (x"ffffffffffffffffffbdef7a039cef39cfdfffffffffffffff"),
                (x"ffffffffffffffffffbdef7a039cef39cfdfffffffffffffff"),
                (x"fffffffffffffffffffdef7a039def7f7bffffffffffffffff"),
                (x"fffffffffffffffffffff8000ef7bde801ffffffffffffffff"),
                (x"fffffffffffffffffffffffffef7ddefffffffffffffffffff"),

                -- 6_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffff4a53bded29def7bda529ffffffffffffffff"),
                (x"ffffffffffa529def874a7bdef7bddef7bda7fffffffffffff"),
                (x"fffffffff4ef7a3f0fbef0c7def7bda529ded3ffffffffffff"),
                (x"fffffffffdf77a31fbc31fbbdf7bdef77bda7694ffffffffff"),
                (x"fffffffffdf77a31fbc31fbbdf7bdef77bda7694ffffffffff"),
                (x"fffffffffd1f7be1f87ef7694a5294efbdded29407ffffffff"),
                (x"fffffffff4f529df769dea6f74a694a529def69407ffffffff"),
                (x"ffffffffffea53ded2f7bdef7bdd3def7b4a5294a03fffffff"),
                (x"ffffffffffea53ded2f7bdef7bdd3def7b4a5294a03fffffff"),
                (x"ffffffffff65ef7bdef7bdef7bdd34a77bdef694a03fffffff"),
                (x"ffffffffff02537bdee94f597bdd34a5294a5294a03fffffff"),
                (x"ffffffffffa3197ba7bded129bdd3de8014a7694003fffffff"),
                (x"fffffffffffd297bf694a3137bdfb4ef7b4a7694003fffffff"),
                (x"fffffffffff8017ba400016f7bde9da77b4a7694a03fffffff"),
                (x"fffffffffff8017ba400016f7bde9da77b4a7694a03fffffff"),
                (x"fffffffffff8017bdc00012f7bde9ea5294ed3bda03fffffff"),
                (x"fffffffffff8017bdf9ce12f7bde9ee8014ed3bda53fffffff"),
                (x"fffffffffff8017bddce712f7bde9ee8000a53bda53fffffff"),
                (x"fffffffffff8017bdef7bdef7bde9ee8000a03bda53fffffff"),
                (x"fffffffffff8017bdef7bdef7bde9ee8000a03bda53fffffff"),
                (x"fffffffffff8009bdef7bdef74a69ea0000003bda53fffffff"),
                (x"fffffffffffffe04def7bdee96319da5280003bda03fffffff"),
                (x"fffffffffffffff0018c6318cf799402520003bda03fffffff"),
                (x"fffffffffffffffff809498d07bcc04def70029407ffffffff"),
                (x"fffffffffffffffff809498d07bcc04def70029407ffffffff"),
                (x"ffffffffffffffff3e1ef40a5f79e94def7f029407ffffffff"),
                (x"fffffffffffffff63fcf7c0b07bde94def748000ffffffffff"),
                (x"fffffffffffffec4f9f08421031bd04def7483ffffffffffff"),
                (x"fffffffffffffe04f9f08421000009bdee9f03ffffffffffff"),
                (x"fffffffffffffe04f9f08421000009bdee9f03ffffffffffff"),
                (x"fffffffffffffff003cf7bdfe4a6f7bdee907fffffffffffff"),
                (x"ffffffffffffffff80c6318c0bdef7ba52c07fffffffffffff"),
                (x"ffffffffffffffffffa73bde04a6e960000fffffffffffffff"),
                (x"ffffffffffffffffffbdef4fd00000ef7a0fffffffffffffff"),
                (x"ffffffffffffffffffbdef4fd00000ef7a0fffffffffffffff"),
                (x"fffffffffffffffffcef7bcfd00000ef7bdfffffffffffffff"),
                (x"ffffffffffffffff83bde9fa00001de8000fffffffffffffff"),
                (x"ffffffffffffffff83c52fba0fffffffffffffffffffffffff")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 3359 := 0;
    signal out_color_reg : std_logic_vector(0 to 199) := (others => '0');
begin
    process(in_sprite_id, in_sprite_row, in_sprite_col, in_sprite_state, in_sprite_direction)
    begin
        real_row <= 0;
        case in_sprite_id is
            when 0 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= in_sprite_row;
                            when D_RIGHT => real_row <= 40 + in_sprite_row;
                            when D_DOWN => real_row <= 80 + in_sprite_row;
                            when D_LEFT => real_row <= 120 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 160 + in_sprite_row;
                            when D_RIGHT => real_row <= 200 + in_sprite_row;
                            when D_DOWN => real_row <= 240 + in_sprite_row;
                            when D_LEFT => real_row <= 280 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 320 + in_sprite_row;
                            when D_RIGHT => real_row <= 360 + in_sprite_row;
                            when D_DOWN => real_row <= 400 + in_sprite_row;
                            when D_LEFT => real_row <= 440 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 1 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 480 + in_sprite_row;
                            when D_RIGHT => real_row <= 520 + in_sprite_row;
                            when D_DOWN => real_row <= 560 + in_sprite_row;
                            when D_LEFT => real_row <= 600 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 640 + in_sprite_row;
                            when D_RIGHT => real_row <= 680 + in_sprite_row;
                            when D_DOWN => real_row <= 720 + in_sprite_row;
                            when D_LEFT => real_row <= 760 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 800 + in_sprite_row;
                            when D_RIGHT => real_row <= 840 + in_sprite_row;
                            when D_DOWN => real_row <= 880 + in_sprite_row;
                            when D_LEFT => real_row <= 920 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 2 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 960 + in_sprite_row;
                            when D_RIGHT => real_row <= 1000 + in_sprite_row;
                            when D_DOWN => real_row <= 1040 + in_sprite_row;
                            when D_LEFT => real_row <= 1080 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1120 + in_sprite_row;
                            when D_RIGHT => real_row <= 1160 + in_sprite_row;
                            when D_DOWN => real_row <= 1200 + in_sprite_row;
                            when D_LEFT => real_row <= 1240 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1280 + in_sprite_row;
                            when D_RIGHT => real_row <= 1320 + in_sprite_row;
                            when D_DOWN => real_row <= 1360 + in_sprite_row;
                            when D_LEFT => real_row <= 1400 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 3 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1440 + in_sprite_row;
                            when D_RIGHT => real_row <= 1480 + in_sprite_row;
                            when D_DOWN => real_row <= 1520 + in_sprite_row;
                            when D_LEFT => real_row <= 1560 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1600 + in_sprite_row;
                            when D_RIGHT => real_row <= 1640 + in_sprite_row;
                            when D_DOWN => real_row <= 1680 + in_sprite_row;
                            when D_LEFT => real_row <= 1720 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1760 + in_sprite_row;
                            when D_RIGHT => real_row <= 1800 + in_sprite_row;
                            when D_DOWN => real_row <= 1840 + in_sprite_row;
                            when D_LEFT => real_row <= 1880 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 4 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1920 + in_sprite_row;
                            when D_RIGHT => real_row <= 1960 + in_sprite_row;
                            when D_DOWN => real_row <= 2000 + in_sprite_row;
                            when D_LEFT => real_row <= 2040 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2080 + in_sprite_row;
                            when D_RIGHT => real_row <= 2120 + in_sprite_row;
                            when D_DOWN => real_row <= 2160 + in_sprite_row;
                            when D_LEFT => real_row <= 2200 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2240 + in_sprite_row;
                            when D_RIGHT => real_row <= 2280 + in_sprite_row;
                            when D_DOWN => real_row <= 2320 + in_sprite_row;
                            when D_LEFT => real_row <= 2360 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 5 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2400 + in_sprite_row;
                            when D_RIGHT => real_row <= 2440 + in_sprite_row;
                            when D_DOWN => real_row <= 2480 + in_sprite_row;
                            when D_LEFT => real_row <= 2520 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2560 + in_sprite_row;
                            when D_RIGHT => real_row <= 2600 + in_sprite_row;
                            when D_DOWN => real_row <= 2640 + in_sprite_row;
                            when D_LEFT => real_row <= 2680 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2720 + in_sprite_row;
                            when D_RIGHT => real_row <= 2760 + in_sprite_row;
                            when D_DOWN => real_row <= 2800 + in_sprite_row;
                            when D_LEFT => real_row <= 2840 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 6 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2880 + in_sprite_row;
                            when D_RIGHT => real_row <= 2920 + in_sprite_row;
                            when D_DOWN => real_row <= 2960 + in_sprite_row;
                            when D_LEFT => real_row <= 3000 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 3040 + in_sprite_row;
                            when D_RIGHT => real_row <= 3080 + in_sprite_row;
                            when D_DOWN => real_row <= 3120 + in_sprite_row;
                            when D_LEFT => real_row <= 3160 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 3200 + in_sprite_row;
                            when D_RIGHT => real_row <= 3240 + in_sprite_row;
                            when D_DOWN => real_row <= 3280 + in_sprite_row;
                            when D_LEFT => real_row <= 3320 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= rom(real_row);
        end if;
    end process;
    out_color <= out_color_reg((in_sprite_col * 5) to ((in_sprite_col + 1) * 5) - 1);
end behavioral;
