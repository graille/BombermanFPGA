library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.PROJECT_PARAMS_PKG.all;
use work.PROJECT_TYPES_PKG.all;
use work.PROJECT_DIRECTION_PKG.all;

entity characters_sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_id : in block_category_type;
        in_sprite_state : in state_type;
        in_sprite_direction : in direction_type;

        in_sprite_row : in integer range 0 to 39;
        in_sprite_col : in integer range 0 to 39;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end characters_sprite_rom;

architecture behavioral of characters_sprite_rom is
    subtype word_t is std_logic_vector(199 downto 0);
    type memory_t is array(3359 downto 0) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- 0_character_0_0
                (x"fffffffffffffffffe94a529def694a53fffffffffffffffff"),
                (x"ffffffffffffff4a53ac677ac633bd67694a5294ffffffffff"),
                (x"ffffffffffffe9def58c1b18c1b18cef58c60d9da53fffffff"),
                (x"ffffffffffffe9def58c1b18c1b18cef58c60d9da53fffffff"),
                (x"fffffffffffd3acef5831b18318d8ceb1831b3b4ffffffffff"),
                (x"fffffffffffd1836318c1b18318fbd6306c677bda53fffffff"),
                (x"ffffffffffa758318d8c1b18c1b18c6319deb0636329ffffff"),
                (x"ffffffffffa758318d8c1b18c1b18c6319deb0636329ffffff"),
                (x"ffffffffffa77ac18d8c6318c1b18c633ac60d9def7b4fffff"),
                (x"ffffffffffa77ac6306c6318c6318c6318c677b4a529ffffff"),
                (x"ffffffffffa77bd6306ceb18ceb18c6319def694a529ffffff"),
                (x"ffffffffffa759d6318ceb18ceb18ceb19def7b4a529ffffff"),
                (x"ffffffffffa758cef59def7acef58ceb194a53bda529ffffff"),
                (x"ffffffffffa758cef59def7acef58ceb194a53bda529ffffff"),
                (x"ffffffffff0518ca53bda77aceb3bda33b4a529d003fffffff"),
                (x"ffffffffff053acef7bda77bdeb3bda77b4a7694003fffffff"),
                (x"fffffffffff829def59def7bdeb3bda53b4a77a0ffffffffff"),
                (x"fffffffffff829da518ceb19da77bded294a7680ffffffffff"),
                (x"fffffffffff829da518ceb19da77bded294a7680ffffffffff"),
                (x"ffffffffffffc14a53aceb9c8bd5ceed294a501fffffffffff"),
                (x"fffffffffffffe0a529dea10ea3ab5ed3b4a53ffffffffffff"),
                (x"ffffffffffff9e4a5294ed6b4ed2b5ed294a11feffffffffff"),
                (x"ffffffffff7902121034eb9dd675cee8004204247bffffffff"),
                (x"ffffffffff7902121034eb9dd675cee8004204247bffffffff"),
                (x"ffffffffff28421294210d28c1b2940842528421297fffffff"),
                (x"fffffffdef094a47bc81277a318e942048f790a5085fffffff"),
                (x"ffffffffde204257bc840d29d1f6940908f79421213dffffff"),
                (x"fffffffd8c4b19e000a10843467694084a00798c4a59ffffff"),
                (x"fffffffd8c4b19e000a10843467694084a00798c4a59ffffff"),
                (x"fffffffc004dd20a53c521094ed084217dde81374a41ffffff"),
                (x"ffffffffff0000ca5294f3df4ebdeff5294a3000003fffffff"),
                (x"fffffffffffffe0a518c6318ca318c63194a03ffffffffffff"),
                (x"fffffffffffffffa518c6318ca318c63194a7fffffffffffff"),
                (x"fffffffffffffffa518c6318ca318c63194a7fffffffffffff"),
                (x"fffffffffffffffa528c63194a518c63294a7fffffffffffff"),
                (x"fffffffffffffff00294a529405294a528007fffffffffffff"),
                (x"fffffffffffffff0029465294052946528007fffffffffffff"),
                (x"fffffffffffffffffc0c63180f818c6301ffffffffffffffff"),
                (x"fffffffffffffffffc0c63180f818c6301ffffffffffffffff"),
                (x"fffffffffffffffffc1df77a0f83bdf741ffffffffffffffff"),

                -- 0_character_0_1
                (x"fffffffffffffffffe94a77bded294ed294a7fffffffffffff"),
                (x"ffffffffffffff4a53ac60c63677bda77bded29fffffffffff"),
                (x"fffffffffffd29d6318318c631b18cef69def7b4ffffffffff"),
                (x"fffffffffffd29d6318318c631b18cef69def7b4ffffffffff"),
                (x"ffffffffffa77ac6319deb18c60d8ced3ac633b4ffffffffff"),
                (x"fffffffffffd29da53ac60c63677bd6758c60d9da53fffffff"),
                (x"fffffffffffd3bdef7b4eb1831b3bda528c60c7da53fffffff"),
                (x"fffffffffffd3bdef7b4eb1831b3bda528c60c7da53fffffff"),
                (x"ffffffffffa77acef7bded28ceb1294a69de8d9da53fffffff"),
                (x"ffffffffffa759def7ac677b44a6f7bdd34a0fbda53fffffff"),
                (x"ffffffffffa759d630631b189bdef7bdef4a33b4ffffffffff"),
                (x"ffffffffffa768c18d8cef7b7bdef7bdefdeb280ffffffffff"),
                (x"ffffffffffa53acef7b4a77b7ba58c632fdef41fffffffffff"),
                (x"ffffffffffa53acef7b4a77b7ba58c632fdef41fffffffffff"),
                (x"ffffffffffa53bda5294ef7b7ba4a5002fded01fffffffffff"),
                (x"fffffffffffd3b4a53b7ef7b7ba484002f4a5c1fffffffffff"),
                (x"fffffffffffd29def697ea537bdc84ef6e94dc1fffffffffff"),
                (x"ffffffffff73bbda5294a2537bdc84f7af7bdc1fffffffffff"),
                (x"ffffffffff73bbda5294a2537bdc84f7af7bdc1fffffffffff"),
                (x"ffffffffff722bd00294a2537bdef7bdef7bdc1fffffffffff"),
                (x"ffffffffbdeb90e00294a3197bdef7bdef7ba41fffffffffff"),
                (x"ffffffd18c675d4ffe94a528cbdef7bdee9483ffffffffffff"),
                (x"ffffffb18ced3fffffc4214be6318c6300007fffffffffffff"),
                (x"ffffffb18ced3fffffc4214be6318c6300007fffffffffffff"),
                (x"ffffffd18ced3fff78810908f2bdef603dffffffffffffffff"),
                (x"ffffffd3bda7ffe295e57bde5f0421630bef7fffffffffffff"),
                (x"ffffffd3bda7ffe7bc81094aff782165bdef7fffffffffffff"),
                (x"ffffffd294ffffe210bef318c003de2b19ef7fffffffffffff"),
                (x"ffffffd294ffffe210bef318c003de2b19ef7fffffffffffff"),
                (x"fffffff7fffffe029597ba537ba4000d99ef7fffffffffffff"),
                (x"fffffffffffffe0632f7bdef7bdc002599ef7fffffffffffff"),
                (x"fffffffffffffff00137ba537ba4002dbdffffffffffffffff"),
                (x"fffffffffffffffffc006318c0018c677fffffffffffffffff"),
                (x"fffffffffffffffffc006318c0018c677fffffffffffffffff"),
                (x"fffffffffffffffffc14a5294a318ca77fffffffffffffffff"),
                (x"ffffffffffffffffffe0a52946318cefffffffffffffffffff"),
                (x"ffffffffffffffffffe0a528c63294ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0528c63000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0528c63000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff077be2f800ffffffffffffffffffff"),

                -- 0_character_0_2
                (x"fffffffffffffffffe94ed29deb294a529ffffffffffffffff"),
                (x"fffffffffffd294a53ac6528c1b3bd677b4a53ffffffffffff"),
                (x"ffffffffffa74636318c677ac1f58c1b3bdef69fffffffffff"),
                (x"ffffffffffa74636318c677ac1f58c1b3bdef69fffffffffff"),
                (x"fffffffffffd3ac18d9def7ac630631b3bdeb3b4ffffffffff"),
                (x"ffffffffffa77bd6306cef7ac6758c677ac60d94ffffffffff"),
                (x"fffffffe9460c6cef59ded28c1f7bded3a318d9da53fffffff"),
                (x"fffffffe9460c6cef59ded28c1f7bded3a318d9da53fffffff"),
                (x"ffffffd18c1b183633b46319d1f7bda329deb3b4a53fffffff"),
                (x"fffffff694a77acef589ba53d1f7bda259def7bda53fffffff"),
                (x"ffffffd294ed29da5137bdefd1f6946253def58ca53fffffff"),
                (x"fffffffe94ef7b4632f7bdefd676944dd2c6519da53fffffff"),
                (x"fffffffe94eb3b44a6f7bdefded129bdee94f7bda53fffffff"),
                (x"fffffffe94eb3b44a6f7bdefded129bdee94f7bda53fffffff"),
                (x"ffffffffffa759dbdd8c65efda26f763197bd3b4ffffffffff"),
                (x"ffffffffff053bdbdca005ef44def7000b7ba689003fffffff"),
                (x"ffffffffff02409bdc8005ee9bdef700097ba417003fffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"ffffffffffffc0cbdc9ef5ef7bdef7f7897bb01fffffffffff"),
                (x"fffffffffffbca04a6f7bdef7bdef7bdee9480afffffffffff"),
                (x"ffffffffff7902563137bdef7bdef7bdd2c614247bffffffff"),
                (x"fffffffdef284242958c4a537bdd294b18529021295fffffff"),
                (x"fffffffdef284242958c4a537bdd294b18529021295fffffff"),
                (x"ffffffbc84215e4294a17b18c6318c784a5291e52108ffffff"),
                (x"fffff797def10af294a40843ef7821090a52bca4f7bc57ffff"),
                (x"fffff7b1294b09e0008f0bdecb31ef0bc800788c4a52c7ffff"),
                (x"fffff626f7ba58000081794a1614a57848000189bdee967fff"),
                (x"fffff626f7ba58000081794a1614a57848000189bdee967fff"),
                (x"fffff626f74deec001e10842cb3021085e0032f74a6e967fff"),
                (x"ffffff81294deeca53cf2108cb308423fd4a32f74a520fffff"),
                (x"fffffffc004dee0a519ef7bde67bdef7994a02f74a41ffffff"),
                (x"ffffffffff0001fa518c6318c6318c63194a7c00003fffffff"),
                (x"ffffffffff0001fa518c6318c6318c63194a7c00003fffffff"),
                (x"fffffffffffffffef68c63194ed18c6329deffffffffffffff"),
                (x"fffffffffffffff0028c631940518c6328007fffffffffffff"),
                (x"fffffffffffffff0028c631940518c6328007fffffffffffff"),
                (x"fffffffffffffffffc14a5280f8294a501ffffffffffffffff"),
                (x"fffffffffffffffffc14a5280f8294a501ffffffffffffffff"),
                (x"ffffffffffffffffffbdf77a0f83bdf77bffffffffffffffff"),

                -- 0_character_0_3
                (x"fffffffffffffffa529def7bdef694a7ffffffffffffffffff"),
                (x"fffffa758c1f694ef5831b18c6318ced29ffffffffffffffff"),
                (x"ffffffd3bd60fac63183677ac1b3bd633b4a7fffffffffffff"),
                (x"ffffffd3bd60fac63183677ac1b3bd633b4a7fffffffffffff"),
                (x"fffffffe94eb3ac6318ceb1836318c18c6c653ffffffffffff"),
                (x"fffffffe94ef7bd6319d60c6c60c631b18c6769fffffffffff"),
                (x"ffffffd3bd633ac18d9deb19d60c63677bdef69fffffffffff"),
                (x"ffffffd3bd633ac18d9deb19d60c63677bdef69fffffffffff"),
                (x"fffffa758cef7a3633b4677bda77bdeb18c6769fffffffffff"),
                (x"ffffffd3bded1836328c4a52cef58c60c631b3b4ffffffffff"),
                (x"fffffffe94a5063ef589bdee9653bdeb18c677b4ffffffffff"),
                (x"ffffffffff0746cef537bdef74d18c677ac677b4ffffffffff"),
                (x"ffffffffff0759d4a58c65ef7bd3bd633b4a769fffffffffff"),
                (x"ffffffffff0759d4a58c65ef7bd3bd633b4a769fffffffffff"),
                (x"fffffffffffd3a9bdc002a537bb294a77bded29fffffffffff"),
                (x"fffffffffff8137bdc0022537bb3bded29def69fffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba694bf7bded01fffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba694a769def5ceffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba694a769def5ceffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694a501ded50effffffffff"),
                (x"fffffffffff8137bdef7bdef7bb294a500e721ddef7fffffff"),
                (x"ffffffffffffc09bdef7bdef765294a03f4a3bac633bffffff"),
                (x"fffffffffffffe00018c6318cf148427bffffe9d6329ffffff"),
                (x"fffffffffffffe00018c6318cf148427bffffe9d6329ffffff"),
                (x"ffffffffffffffff780c7bde579021093dfffe9d6329ffffff"),
                (x"ffffffffffffffe2958c0843e2bdef2bcbef7ff4ef69ffffff"),
                (x"ffffffffffffffef7acc0fbde79421091fef7fffef69ffffff"),
                (x"ffffffffffffffe63185f0000633def149ef7ffffffbffffff"),
                (x"ffffffffffffffe63185f0000633def149ef7ffffffbffffff"),
                (x"ffffffffffffffe632c102537ba6f7bb0a007fffffffffffff"),
                (x"ffffffffffffffe632c405ef7bdef7bdd8007fffffffffffff"),
                (x"ffffffffffffffff7ac502537ba6f7ba41ffffffffffffffff"),
                (x"ffffffffffffffffffac600006318c003fffffffffffffffff"),
                (x"ffffffffffffffffffac600006318c003fffffffffffffffff"),
                (x"ffffffffffffffffffb463194a5294a03fffffffffffffffff"),
                (x"fffffffffffffffffffd6318ca529407ffffffffffffffffff"),
                (x"ffffffffffffffffffffa318c6529407ffffffffffffffffff"),
                (x"ffffffffffffffffffff0318c65000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0318c65000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc5f7400ffffffffffffffffffff"),

                -- 0_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a529def694a53fffffffffffffffff"),
                (x"ffffffffffffff4a53ac677ac633bd67694a5294ffffffffff"),
                (x"ffffffffffffff4a53ac677ac633bd67694a5294ffffffffff"),
                (x"ffffffffffffe9def58c1b18c1b18cef58c60d9da53fffffff"),
                (x"fffffffffffd3acef5831b18318d8ceb1831b3b4ffffffffff"),
                (x"fffffffffffd1836318c1b18318fbd6306c677bda53fffffff"),
                (x"fffffffffffd1836318c1b18318fbd6306c677bda53fffffff"),
                (x"ffffffffffa758318d8c1b18c1b18c6319deb0636329ffffff"),
                (x"ffffffffffa77ac18d8c6318c1b18c633ac60d9def7b4fffff"),
                (x"ffffffffffa77ac6306c6318c6318c6318c677b4a529ffffff"),
                (x"ffffffffffa77bd6306ceb18ceb18c6319def694a529ffffff"),
                (x"ffffffffffa759d6318ceb18ceb18ceb19def7b4a529ffffff"),
                (x"ffffffffffa759d6318ceb18ceb18ceb19def7b4a529ffffff"),
                (x"ffffffffffa758cef59def7acef58ceb194a53bda529ffffff"),
                (x"ffffffffff0518ca53bda77aceb3bda33b4a529d003fffffff"),
                (x"ffffffffff053acef7bda77bdeb3bda77b4a7694003fffffff"),
                (x"fffffffffff829def59def7bdeb3bda53b4a77a0ffffffffff"),
                (x"fffffffffff829def59def7bdeb3bda53b4a77a0ffffffffff"),
                (x"fffffffffff829da518ceb19da77bded294a7680ffffffffff"),
                (x"ffffffffffffc14a53aceb9c8bd5ceed294a501fffffffffff"),
                (x"fffffffffffffc0a529dea10ea3ab5ed3b4a53ffffffffffff"),
                (x"ffffffffffff8a4a5294ed6b4ed2b5ed294a13dfffffffffff"),
                (x"ffffffffffff8a4a5294ed6b4ed2b5ed294a13dfffffffffff"),
                (x"fffffffffff148429434eb9dd633bde80010849effffffffff"),
                (x"fffffffffff10a57bc210d28c18d8c090a10843effffffffff"),
                (x"fffffffffff1484f78240f7ac18d8c090a108485f7bfffffff"),
                (x"ffffffffff67bde7bc810843460fbd091e529484f7bfffffff"),
                (x"ffffffffff67bde7bc810843460fbd091e529484f7bfffffff"),
                (x"ffffffffff031807bca408421eb294295e10843e633fffffff"),
                (x"fffffffffff8000f79e529084a7694f781ef7bc9633fffffff"),
                (x"fffffffffffffffef69463194a5294a53ac62520ffffffffff"),
                (x"fffffffffffffffef6946318ca518c653bde801fffffffffff"),
                (x"fffffffffffffffef6946318ca518c653bde801fffffffffff"),
                (x"fffffffffffffffef7b4a318ca77bdef40007fffffffffffff"),
                (x"fffffffffffffffffc1da529460294a03fffffffffffffffff"),
                (x"ffffffffffffffffffe0eb18ce800007ffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc3f03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc3f03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bdde83ffffffffffffffffffffff"),

                -- 0_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bded294ed294a7fffffffffffff"),
                (x"ffffffffffffff4a53ac60c63677bda77bded29fffffffffff"),
                (x"ffffffffffffff4a53ac60c63677bda77bded29fffffffffff"),
                (x"fffffffffffd29d6318318c631b18cef69def7b4ffffffffff"),
                (x"ffffffffffa77ac6319deb18c60d8ced3ac633b4ffffffffff"),
                (x"fffffffffffd29da53ac60c63677bd6758c60d9da53fffffff"),
                (x"fffffffffffd29da53ac60c63677bd6758c60d9da53fffffff"),
                (x"fffffffffffd3bdef7b4eb1831b3bda528c60c7da53fffffff"),
                (x"ffffffffffa77acef7bded28ceb1294a69de8d9da53fffffff"),
                (x"ffffffffffa759def7ac677b44a6f7bdd34a0fbda53fffffff"),
                (x"ffffffffffa759d630631b189bdef7bdef4a33b4ffffffffff"),
                (x"ffffffffffa768c18d8cef7b7bdef7bdefdeb280ffffffffff"),
                (x"ffffffffffa768c18d8cef7b7bdef7bdefdeb280ffffffffff"),
                (x"ffffffffffa53acef7b4a77b7ba58c632fdef41fffffffffff"),
                (x"ffffffffffa53bda5294ef7b7ba4a5002fded01fffffffffff"),
                (x"fffffffffffd3b4a53b7ef7b7ba484002f4a5c1fffffffffff"),
                (x"fffffffffffd29def697ea537bdc84ef6e94dc1fffffffffff"),
                (x"fffffffffffd29def697ea537bdc84ef6e94dc1fffffffffff"),
                (x"ffffffffff73bbda5294a2537bdc84f7af7bdc1fffffffffff"),
                (x"ffffffffff722bd00294a2537bdef7bdef7bdc1fffffffffff"),
                (x"fffffffe94eb90e00294a3197bdef7bdef7ba41fffffffffff"),
                (x"fffffff58c675d4ffe94a528cbdef7bdee9483ffffffffffff"),
                (x"fffffff58c675d4ffe94a528cbdef7bdee9483ffffffffffff"),
                (x"ffffffd18ced3ff003c5214af6318c6300007fffffffffffff"),
                (x"ffffffd3bda7fff000a408425f3def783dffffffffffffffff"),
                (x"ffffffd294fffe0f7884294a47f8842798007fffffffffffff"),
                (x"ffffffd3fffffe0f78af08421f17de2798007fffffffffffff"),
                (x"ffffffd3fffffe0f78af08421f17de2798007fffffffffffff"),
                (x"fffffffffffffe07bde42bdfef000003cac67fffffffffffff"),
                (x"fffffffffffffe07bfc5f318965ef7b80ac67fffffffffffff"),
                (x"fffffffffffffe0f79e04def74def7b81ec67fffffffffffff"),
                (x"ffffffffffffff4003de025374a6f76501ffffffffffffffff"),
                (x"ffffffffffffff4003de025374a6f76501ffffffffffffffff"),
                (x"ffffffffffffff4a518ca000c60000053fffffffffffffffff"),
                (x"fffffffffffffe0a518c6529405294a7ffffffffffffffffff"),
                (x"fffffffffffffe0a528ca52940518c653fffffffffffffffff"),
                (x"fffffffffffffff0018c6528000294f7bfffffffffffffffff"),
                (x"fffffffffffffff0018c6528000294f7bfffffffffffffffff"),
                (x"fffffffffffffff003be2fbc0fffffffffffffffffffffffff"),

                -- 0_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ed29deb294a529ffffffffffffffff"),
                (x"fffffffffffd294a53ac6528c1b3bd677b4a53ffffffffffff"),
                (x"fffffffffffd294a53ac6528c1b3bd677b4a53ffffffffffff"),
                (x"ffffffffffa74636318c677ac1f58c1b3bdef69fffffffffff"),
                (x"fffffffffffd3ac18d9def7ac630631b3bdeb3b4ffffffffff"),
                (x"ffffffffffa77bd6306cef7ac6758c677ac60d94ffffffffff"),
                (x"ffffffffffa77bd6306cef7ac6758c677ac60d94ffffffffff"),
                (x"fffffffe9460c6cef59ded28c1f7bded3a318d9da53fffffff"),
                (x"ffffffd18c1b183633b46319d1f7bda329deb3b4a53fffffff"),
                (x"fffffff694a77acef589ba53d1f7bda259def7bda53fffffff"),
                (x"ffffffd294ed29da5137bdefd1f6946253def58ca53fffffff"),
                (x"fffffffe94ef7b4632f7bdefd676944dd2c6519da53fffffff"),
                (x"fffffffe94ef7b4632f7bdefd676944dd2c6519da53fffffff"),
                (x"fffffffe94eb3b44a6f7bdefded129bdee94f7bda53fffffff"),
                (x"ffffffffffa759dbdd8c65efda26f763197bd3b4ffffffffff"),
                (x"ffffffffff053bdbdca005ef44def7000b7ba689003fffffff"),
                (x"ffffffffff02409bdc8005ee9bdef700097ba417003fffffff"),
                (x"ffffffffff02409bdc8005ee9bdef700097ba417003fffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"ffffffffffffc0cbdc9ef5ef7bdef7f7897bb01fffffffffff"),
                (x"ffffffffffff9e04a6f7bdef7bdef7bdee9483deffffffffff"),
                (x"ffffffffff7948563137bdef7bdef7bdd2c61424f7bfffffff"),
                (x"ffffffffff7948563137bdef7bdef7bdd2c61424f7bfffffff"),
                (x"fffffffdef290842958c4a537bdd294b18f78484297dffffff"),
                (x"fffffff88423ca4211e17b18c6318c791e52bc21210befffff"),
                (x"fffffff9ef291ef295e40843ef7821091ef791ef7bcbefffff"),
                (x"ffffffb12963ca07bc8f0bdecb31ef0bc8f78129633dffffff"),
                (x"ffffffb12963ca07bc8f0bdecb31ef0bc8f78129633dffffff"),
                (x"ffffffb1294b1807bc81794a1614a578400032f74a59ffffff"),
                (x"ffffffb2f7ba41f7bca10842cb302109597bdee94a59ffffff"),
                (x"ffffffb129bb01fa53de2908cb30a5f7997bdd2c6301ffffff"),
                (x"ffffff81294b3ffa518c6318c6318c650094dd80003fffffff"),
                (x"ffffff81294b3ffa518c6318c6318c650094dd80003fffffff"),
                (x"fffffffc00003ffa528c6318ca5294a52800001fffffffffff"),
                (x"fffffffffffffffffe8c6318c60294a529ffffffffffffffff"),
                (x"fffffffffffffffffff46318c603bdef7fffffffffffffffff"),
                (x"ffffffffffffffffffe0a529de800007ffffffffffffffffff"),
                (x"ffffffffffffffffffe0a529de800007ffffffffffffffffff"),
                (x"ffffffffffffffffffffef7beeffffffffffffffffffffffff"),

                -- 0_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa529def7bdef694a7ffffffffffffffffff"),
                (x"fffffa758c1f694ef5831b18c6318ced29ffffffffffffffff"),
                (x"fffffa758c1f694ef5831b18c6318ced29ffffffffffffffff"),
                (x"ffffffd3bd60fac63183677ac1b3bd633b4a7fffffffffffff"),
                (x"fffffffe94eb3ac6318ceb1836318c18c6c653ffffffffffff"),
                (x"fffffffe94ef7bd6319d60c6c60c631b18c6769fffffffffff"),
                (x"fffffffe94ef7bd6319d60c6c60c631b18c6769fffffffffff"),
                (x"ffffffd3bd633ac18d9deb19d60c63677bdef69fffffffffff"),
                (x"fffffa758cef7a3633b4677bda77bdeb18c6769fffffffffff"),
                (x"ffffffd3bded1836328c4a52cef58c60c631b3b4ffffffffff"),
                (x"fffffffe94a5063ef589bdee9653bdeb18c677b4ffffffffff"),
                (x"ffffffffff0746cef537bdef74d18c677ac677b4ffffffffff"),
                (x"ffffffffff0746cef537bdef74d18c677ac677b4ffffffffff"),
                (x"ffffffffff0759d4a58c65ef7bd3bd633b4a769fffffffffff"),
                (x"fffffffffffd189bdc002a537bb294a77bded29fffffffffff"),
                (x"fffffffffff8137bdc0022537bb3bded29def69fffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba694bf7bded01fffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba694bf7bded01fffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba694a769def5ceffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694a501ded50effffffffff"),
                (x"fffffffffff8137bdef7bdef7bb294a500e721dda53fffffff"),
                (x"ffffffffffffc09bdef7bdef765294a03f4a3bac633bffffff"),
                (x"ffffffffffffc09bdef7bdef765294a03f4a3bac633bffffff"),
                (x"fffffffffffffe00018c6318c794842f81fffe9d6329ffffff"),
                (x"ffffffffffffffff780f7bdfe284212141fffff4ef69ffffff"),
                (x"fffffffffffffe0633c427bcf214a5213c007fffa529ffffff"),
                (x"fffffffffffffe0633c4f14be08421797c007fffffe9ffffff"),
                (x"fffffffffffffe0633c4f14be08421797c007fffffe9ffffff"),
                (x"fffffffffffffec295e00001ef3ca523de007fffffffffffff"),
                (x"fffffffffffffec29417bdeec4b3de2f9e007fffffffffffff"),
                (x"fffffffffffffec7bc17bdee9bdd2903fc007fffffffffffff"),
                (x"fffffffffffffff0028cba529ba400f7814a7fffffffffffff"),
                (x"fffffffffffffff0028cba529ba400f7814a7fffffffffffff"),
                (x"fffffffffffffffffe800000c6029463294a7fffffffffffff"),
                (x"fffffffffffffffffff4a5280a518c6328007fffffffffffff"),
                (x"fffffffffffffffffe8c65280a52946528007fffffffffffff"),
                (x"ffffffffffffffffffdea00000518c6301ffffffffffffffff"),
                (x"ffffffffffffffffffdea00000518c6301ffffffffffffffff"),
                (x"fffffffffffffffffffffffff078a5f741ffffffffffffffff"),

                -- 0_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a529def694a53fffffffffffffffff"),
                (x"ffffffffffffff4a53ac677ac633bd67694a5294ffffffffff"),
                (x"ffffffffffffff4a53ac677ac633bd67694a5294ffffffffff"),
                (x"ffffffffffffe9def58c1b18c1b18cef58c60d9da53fffffff"),
                (x"fffffffffffd3acef5831b18318d8ceb1831b3b4ffffffffff"),
                (x"fffffffffffd1836318c1b18318fbd6306c677bda53fffffff"),
                (x"fffffffffffd1836318c1b18318fbd6306c677bda53fffffff"),
                (x"ffffffffffa758318d8c1b18c1b18c6319deb0636329ffffff"),
                (x"ffffffffffa77ac18d8c6318c1b18c633ac60d9def7b4fffff"),
                (x"ffffffffffa77ac6306c6318c6318c6318c677b4a529ffffff"),
                (x"ffffffffffa77bd6306ceb18ceb18c6319def694a529ffffff"),
                (x"ffffffffffa759d6318ceb18ceb18ceb19def7b4a529ffffff"),
                (x"ffffffffffa759d6318ceb18ceb18ceb19def7b4a529ffffff"),
                (x"ffffffffffa758cef59def7acef58ceb194a53bda529ffffff"),
                (x"ffffffffff0518ca53bda77aceb3bda33b4a529d003fffffff"),
                (x"ffffffffff053acef7bda77bdeb3bda77b4a7694003fffffff"),
                (x"fffffffffff829def59def7bdeb3bda53b4a77a0ffffffffff"),
                (x"fffffffffff829def59def7bdeb3bda53b4a77a0ffffffffff"),
                (x"fffffffffff829da518ceb19da77bded294a7680ffffffffff"),
                (x"ffffffffffffc14a53aceb9c8bd5ceed294a501fffffffffff"),
                (x"fffffffffffffe0a529dea10ea3ab5ed3b4a53dfffffffffff"),
                (x"fffffffffffffc4a5294ed6b4ed2b5ed294a10beffffffffff"),
                (x"fffffffffffffc4a5294ed6b4ed2b5ed294a10beffffffffff"),
                (x"ffffffffffff88108494ed29d675cee800529085f7bfffffff"),
                (x"ffffffffffff821084a40f7ac1f6940842f794a4f7bfffffff"),
                (x"fffffffffff1481084a40b1831f6940903ef1085f7bfffffff"),
                (x"fffffffffff1085295e40b183650210848f7fbde633fffffff"),
                (x"fffffffffff1085295e40b183650210848f7fbde633fffffff"),
                (x"ffffffffff67821085e52f7a3ed021090af7818c003fffffff"),
                (x"ffffffffff627def781ef528ca1084295fef0000ffffffffff"),
                (x"fffffffffff8129633b4a529da53bded29deffffffffffffff"),
                (x"ffffffffffffc00ef7b463194a318c6529deffffffffffffff"),
                (x"ffffffffffffc00ef7b463194a318c6529deffffffffffffff"),
                (x"fffffffffffffff0001def7bda318ca53bdeffffffffffffff"),
                (x"ffffffffffffffffffe0a528065294a741ffffffffffffffff"),
                (x"ffffffffffffffffffff00000eb18ce83fffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f0fde07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f0fde07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0ef7de07ffffffffffffffffff"),

                -- 0_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a77bded294ed294a7fffffffffffff"),
                (x"ffffffffffffff4a53ac60c63677bda77bded29fffffffffff"),
                (x"ffffffffffffff4a53ac60c63677bda77bded29fffffffffff"),
                (x"fffffffffffd29d6318318c631b18cef69def7b4ffffffffff"),
                (x"ffffffffffa77ac6319deb18c60d8ced3ac633b4ffffffffff"),
                (x"fffffffffffd29da53ac60c63677bd6758c60d9da53fffffff"),
                (x"fffffffffffd29da53ac60c63677bd6758c60d9da53fffffff"),
                (x"fffffffffffd3bdef7b4eb1831b3bda528c60c7da53fffffff"),
                (x"ffffffffffa77acef7bded28ceb1294a69de8d9da53fffffff"),
                (x"ffffffffffa759def7ac677b44a6f7bdd34a0fbda53fffffff"),
                (x"ffffffffffa759d630631b189bdef7bdef4a33b4ffffffffff"),
                (x"ffffffffffa768c18d8cef7b7bdef7bdefdeb280ffffffffff"),
                (x"ffffffffffa768c18d8cef7b7bdef7bdefdeb280ffffffffff"),
                (x"ffffffffffa53acef7b4a3197ba58c632fdef41fffffffffff"),
                (x"ffffffffffa53bda529463197ba4a5002fded01fffffffffff"),
                (x"fffffffffffd3b4a53b763197ba484002f4a5c1fffffffffff"),
                (x"fffffffffffd29def69762537bdc84ef6e94dc1fffffffffff"),
                (x"fffffffffffd29def69762537bdc84ef6e94dc1fffffffffff"),
                (x"ffffffffff73bbda5294a2537bdc84f7af7bdc1fffffffffff"),
                (x"ffffffffff722bda5294a2537bdef7bdef7bdc1fffffffffff"),
                (x"fffffffe94eb90ea5294a3197bdef7bdef7ba41fffffffffff"),
                (x"fffffffe94675d4a5294a528cbdef7bdee9483ffffffffffff"),
                (x"fffffffe94675d4a5294a528cbdef7bdee9483ffffffffffff"),
                (x"fffffffe946769f000a42fbde6318c6300007fffffffffffff"),
                (x"fffffffe94ed3e02942123de523def483dffffffffffffffff"),
                (x"fffffffe94ed3fe7bc84094be08484610bef7fffffffffffff"),
                (x"fffffffe94a7c0f21021294a57858cb78ac67fffffffffffff"),
                (x"fffffffe94a7c0f21021294a57858cb78ac67fffffffffffff"),
                (x"ffffffffbda7c05f79ef27bcf2798c617c94b3ffffffffffff"),
                (x"ffffffffffa7c1e4a6f7480002118cb17c9483ffffffffffff"),
                (x"fffffffffffffe04a6f7bdee9f158cb780007fffffffffffff"),
                (x"fffffffffffffe063137bdef70318cb501ffffffffffffffff"),
                (x"fffffffffffffe063137bdef70318cb501ffffffffffffffff"),
                (x"fffffffffffffff0000c4dee90318c653fffffffffffffffff"),
                (x"fffffffffffffff0029400000a3294a53fffffffffffffffff"),
                (x"fffffffffffffffef7b400000a318c633fffffffffffffffff"),
                (x"fffffffffffffff0001de80000518cef41ffffffffffffffff"),
                (x"fffffffffffffff0001de80000518cef41ffffffffffffffff"),
                (x"fffffffffffffffffffffffff077de2f81ffffffffffffffff"),

                -- 0_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ed29deb294a529ffffffffffffffff"),
                (x"fffffffffffd294a53ac6528c1b3bd677b4a53ffffffffffff"),
                (x"fffffffffffd294a53ac6528c1b3bd677b4a53ffffffffffff"),
                (x"ffffffffffa74636318c677ac1f58c1b3bdef69fffffffffff"),
                (x"fffffffffffd3ac18d9def7ac630631b3bdeb3b4ffffffffff"),
                (x"ffffffffffa77bd6306cef7ac6758c677ac60d94ffffffffff"),
                (x"ffffffffffa77bd6306cef7ac6758c677ac60d94ffffffffff"),
                (x"fffffffe9460c6cef59ded28c1f7bded3a318d9da53fffffff"),
                (x"ffffffd18c1b183633b46319d1f7bda329deb3b4a53fffffff"),
                (x"fffffff694a77acef589ba53d1f7bda259def7bda53fffffff"),
                (x"ffffffd294ed29da5137bdefd1f6946253def58ca53fffffff"),
                (x"fffffffe94ef7b4632f7bdefd676944dd2c6519da53fffffff"),
                (x"fffffffe94ef7b4632f7bdefd676944dd2c6519da53fffffff"),
                (x"fffffffe94eb3b44a6f7bdefded129bdee94f7bda53fffffff"),
                (x"ffffffffffa759dbdd8c65efda26f763197bd3b4ffffffffff"),
                (x"ffffffffff053bdbdca005ef44def7000b7ba689003fffffff"),
                (x"ffffffffff02409bdc8005ee9bdef700097ba417003fffffff"),
                (x"ffffffffff02409bdc8005ee9bdef700097ba417003fffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"ffffffffffffc0cbdc9ef5ef7bdef7f7897bb01fffffffffff"),
                (x"ffffffffffffbc04a6f7bdef7bdef7bdee9481feffffffffff"),
                (x"fffffffffff102563137bdef7bdef7bdd2c614857bffffffff"),
                (x"fffffffffff102563137bdef7bdef7bdd2c614857bffffffff"),
                (x"ffffffffde290817bd8c4a537bdd294b18529084295fffffff"),
                (x"fffffff8a52042f295e47b18c6318c785e4210af2109efffff"),
                (x"fffffff8a57bde47bde40843ef7821091e52bde4295fefffff"),
                (x"ffffffffde625207bc8f0bdecb31ef0bc8f780af6312cfffff"),
                (x"ffffffffde625207bc8f0bdecb31ef0bc8f780af6312cfffff"),
                (x"fffffffd8c4deec00001794a1614a57848f7818c4a52cfffff"),
                (x"fffffffd8c4a6f7bdd850842cb3021084af7fc09bdeecfffff"),
                (x"fffffffc0063137bdd9ef14acb30842fbd4a7c0cbdd2cfffff"),
                (x"ffffffffff001974a4146318c6318c63194a7fec4a520fffff"),
                (x"ffffffffff001974a4146318c6318c63194a7fec4a520fffff"),
                (x"ffffffffffffc0000294a5294a318c63294a7fe00001ffffff"),
                (x"fffffffffffffffffe94a52806318c6329ffffffffffffffff"),
                (x"fffffffffffffffffffdef7a06318c653fffffffffffffffff"),
                (x"ffffffffffffffffffff00000ef694a03fffffffffffffffff"),
                (x"ffffffffffffffffffff00000ef694a03fffffffffffffffff"),
                (x"fffffffffffffffffffffffffefbbdefffffffffffffffffff"),

                -- 0_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa529def7bdef694a7ffffffffffffffffff"),
                (x"fffffa758c1f694ef5831b18c6318ced29ffffffffffffffff"),
                (x"fffffa758c1f694ef5831b18c6318ced29ffffffffffffffff"),
                (x"ffffffd3bd60fac63183677ac1b3bd633b4a7fffffffffffff"),
                (x"fffffffe94eb3ac6318ceb1836318c18c6c653ffffffffffff"),
                (x"fffffffe94ef7bd6319d60c6c60c631b18c6769fffffffffff"),
                (x"fffffffe94ef7bd6319d60c6c60c631b18c6769fffffffffff"),
                (x"ffffffd3bd633ac18d9deb19d60c63677bdef69fffffffffff"),
                (x"fffffa758cef7a3633b4677bda77bdeb18c6769fffffffffff"),
                (x"ffffffd3bded1836328c4a52cef58c60c631b3b4ffffffffff"),
                (x"fffffffe94a5063ef589bdee9653bdeb18c677b4ffffffffff"),
                (x"ffffffffff0746cef537bdef74d18c677ac677b4ffffffffff"),
                (x"ffffffffff0746cef537bdef74d18c677ac677b4ffffffffff"),
                (x"ffffffffff0759d4a58c65ef7bd3bd633b4a769fffffffffff"),
                (x"fffffffffffd3a9bdc002a537bb294a77bded29fffffffffff"),
                (x"fffffffffff8137bdc0022537bb3bded29def69fffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba694bf7bded01fffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba694bf7bded01fffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba694a769def5ceffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694a501ded50effffffffff"),
                (x"fffffffffff8137bdef7bdef7bb294a528e721ddffffffffff"),
                (x"ffffffffffffc09bdef7bdef765294a0294a3bacef7fffffff"),
                (x"ffffffffffffc09bdef7bdef765294a0294a3bacef7fffffff"),
                (x"fffffffffffffe00018c6318cf78a52141ffd3aca53fffffff"),
                (x"ffffffffffffffff78097bde42bc84084a007e9da53fffffff"),
                (x"ffffffffffffffe2948c20421f1421211fef7e9da53fffffff"),
                (x"fffffffffffffec297d66042f294a50848f783f4a53fffffff"),
                (x"fffffffffffffec297d66042f294a50848f783f4a53fffffff"),
                (x"ffffffffffffd89f78ac67bc47f8847bfc5283ffef7fffffff"),
                (x"ffffffffffffc09f78b66108400129bdd3ef03ffffffffffff"),
                (x"fffffffffffffe0003d6614be4def7bdd2007fffffffffffff"),
                (x"fffffffffffffff0029663180bdef7ba58007fffffffffffff"),
                (x"fffffffffffffff0029663180bdef7ba58007fffffffffffff"),
                (x"fffffffffffffffffe8c631804dd296001ffffffffffffffff"),
                (x"fffffffffffffffffe94a319400000a501ffffffffffffffff"),
                (x"fffffffffffffffffd8c6319400000a77bffffffffffffffff"),
                (x"fffffffffffffff003bd65280003bde801ffffffffffffffff"),
                (x"fffffffffffffff003bd65280003bde801ffffffffffffffff"),
                (x"fffffffffffffff003c5f77a0fffffffffffffffffffffffff"),

                -- 1_character_0_0
                (x"fffffffffffffffef7ae739ddeb9ce73bbdeffffffffffffff"),
                (x"fffffffffffffbd73ab5ab9ce756b5ad6ae73bbdffffffffff"),
                (x"ffffffffffff5d5ad517456aead6b5422e8456aeef7fffffff"),
                (x"ffffffffffff5d5ad517456aead6b5422e8456aeef7fffffff"),
                (x"fffffffffffffae73aa84210eab9ceaa115abbbdffffffffff"),
                (x"ffffffffffff5d5bdd15ab9ce756b575517ba2aeef7fffffff"),
                (x"ffffffffbdebaa8ad6b5ad6b5722b5ab915ad6b573bbffffff"),
                (x"ffffffffbdebaa8ad6b5ad6b5722b5ab915ad6b573bbffffff"),
                (x"fffffff5cead6b5739d5456b572108abaa843ab5ad5ddfffff"),
                (x"ffffffffbd756ae73ab7456ae75ef7ab9d5aa1ddef7bffffff"),
                (x"ffffffffffebab573aa8ad6b5ad508755ce756ae73bfffffff"),
                (x"ffffffffbd756aead6b5aa115756b5756ae73ab573bbffffff"),
                (x"fffffff5ceabbaead6aeaa115755ce73aae739ce739dffffff"),
                (x"fffffff5ceabbaead6aeaa115755ce73aae739ce739dffffff"),
                (x"fffffef7bdef5cead5dd456aeeb9ceef5ce777bd73bbdfffff"),
                (x"ffffffffff076ae73bae456bdebbbd777ae73bbd003fffffff"),
                (x"ffffffffff076aeef7aeab9dd777bd73bae7381d003fffffff"),
                (x"fffffffffff81dd73abd777aeaf5ceabbae77400ffffffffff"),
                (x"fffffffffff81dd73abd777aeaf5ceabbae77400ffffffffff"),
                (x"ffffffffffffc1d73abdeb9ceabab5ab9ddef41fffffffffff"),
                (x"fffffffffffffe0ef5ddeb9d5739ceabbbde83ffffffffffff"),
                (x"fffffffffffffde003aeef7aeef5ce73ba007bdfffffffffff"),
                (x"ffffffffffff8a421000ef7bd077bd70004211feffffffffff"),
                (x"ffffffffffff8a421000ef7bd077bd70004211feffffffffff"),
                (x"fffffffffff14210842500000000000142108425f7bfffffff"),
                (x"fffffffffff042129421294a5294a52842528421f7bfffffff"),
                (x"ffffffffde28421f78a10842108421084bef0421297dffffff"),
                (x"ffffffffde29425000a10842108421084a001425297dffffff"),
                (x"ffffffffde29425000a10842108421084a001425297dffffff"),
                (x"ffffffffdef14a0f78a10842108421084bef00a5f7bdffffff"),
                (x"ffffffffff0001e294210842128421084252f800003fffffff"),
                (x"fffffffffffffe02942108421f042108425283ffffffffffff"),
                (x"ffffffffffffffff78a108425f1421084a217fffffffffffff"),
                (x"ffffffffffffffff78a108425f1421084a217fffffffffffff"),
                (x"ffffffffffffffff7bdef7bdef7bde1084217fffffffffffff"),
                (x"fffffffffffffff00047108420084211c4007fffffffffffff"),
                (x"fffffffffffffff0004739ce2008e739c4007fffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc1425280f82942501ffffffffffffffff"),

                -- 1_character_0_1
                (x"fffffffffffffffffffdef7bdef7bd739ddef7ffffffffffff"),
                (x"ffffffffffffffdef5cead6b5ab9ce75508455ce73bfffffff"),
                (x"ffffffffffff7aead6a8bdef7456b5721084211573bbffffff"),
                (x"ffffffffffff7aead6a8bdef7456b5721084211573bbffffff"),
                (x"ffffffffffeb9d5ad508456b5ad6b5ad6b5ab9ddef7fffffff"),
                (x"ffffffffffff7aead6b5adef7455ce73ab5ad5ddffffffffff"),
                (x"ffffffffffeb9d5ad6a84211573ab5ad5c8422aeef7fffffff"),
                (x"ffffffffffeb9d5ad6a84211573ab5ad5c8422aeef7fffffff"),
                (x"ffffffffffebab5ad508ad6ae756b5457b5adeee73bbffffff"),
                (x"ffffffffbd756b573ab5739ce75508bbbae72115739ddfffff"),
                (x"fffffff5cead5cead6aeeb9ddaa1087759ded515ef7fffffff"),
                (x"ffffffffbdebbb5ad5dd739dd455ceef53debaaeef7fffffff"),
                (x"ffffffffffef6ae73bae777b5abbbd6312c676bdffffffffff"),
                (x"ffffffffffef6ae73bae777b5abbbd6312c676bdffffffffff"),
                (x"ffffffffffeb9ddef7aeeb9d5738a5002e94f5ddffffffffff"),
                (x"ffffffffffef7bdef7bdeb9ceea484002f7ba7bfffffffffff"),
                (x"ffffffffffef7bdef689ef7a9bdc84802f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7b4a2537bdc84842f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7b4a2537bdc84842f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7bda2537bdef7bdef7bdc1fffffffffff"),
                (x"fffffffffffffbf003bda3197bdef7bdef7ba41fffffffffff"),
                (x"fffffffffffffffffe9da528cbdef7bdee9483ffffffffffff"),
                (x"ffffffffffffffffffcf7bde26318c6300007fffffffffffff"),
                (x"ffffffffffffffffffcf7bde26318c6300007fffffffffffff"),
                (x"ffffffffffffffff78a1094a52fa94a53fffffffffffffffff"),
                (x"ffffffffffffffff782108425096941dbdffffffffffffffff"),
                (x"ffffffffffffffe29421294bef14a51b19ffffffffffffffff"),
                (x"ffffffffffffffe084250843e278a5a52dffffffffffffffff"),
                (x"ffffffffffffffe084250843e278a5a52dffffffffffffffff"),
                (x"ffffffffffffffe08421094a44dd8c292dffffffffffffffff"),
                (x"fffffffffffffe0294210fbc34dd8c0d19ffffffffffffffff"),
                (x"fffffffffffffff000a52fbcf62400097dffffffffffffffff"),
                (x"ffffffffffffffff7800f7bde01421097dffffffffffffffff"),
                (x"ffffffffffffffff7800f7bde01421097dffffffffffffffff"),
                (x"fffffffffffffff10bc5294a5084212fbfffffffffffffffff"),
                (x"fffffffffffffffffc42f7bdef7bdef7ffffffffffffffffff"),
                (x"ffffffffffffffffffe011ce739c00ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0084738800ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0084738800ffffffffffffffffffff"),
                (x"ffffffffffffffffffffa529425000ffffffffffffffffffff"),

                -- 1_character_0_2
                (x"fffffffffffffffef7ae739ceef5ce73bbdeffffffffffffff"),
                (x"ffffffffffff7ae73ab5ad6b5739cead6ae777bfffffffffff"),
                (x"ffffffffffebab5422e8456b5abab545d15ad5ddffffffffff"),
                (x"ffffffffffebab5422e8456b5abab545d15ad5ddffffffffff"),
                (x"ffffffffffff7aead508ab9ceab908422ae73bbfffffffffff"),
                (x"ffffffffffebaa8bdd15756b5777bd75517bd5ddffffffffff"),
                (x"ffffffffbd756b5ad50ead6a8775ceabab5aa2aeef7bffffff"),
                (x"ffffffffbd756b5ad50ead6a8775ceabab5aa2aeef7bffffff"),
                (x"fffffff5cead6ae422ae42108777bd455ce756b5ad5ddfffff"),
                (x"ffffffffbdef5c8ad6ae45ef7777bd45dce73ab573bbffffff"),
                (x"ffffffffff73ab573aaeaa115733bd722bdeb9d5ef7fffffff"),
                (x"ffffffffbd756aead6ae756b57258ced6ae775ce73bbffffff"),
                (x"fffffffdceab9cead5ddeb9d5edd29ebaae775ce739ddfffff"),
                (x"fffffffdceab9cead5ddeb9d5edd29ebaae775ce739ddfffff"),
                (x"fffffff7bd777ae73bac677aeedef7675d5af5ddef7bdeffff"),
                (x"ffffffffff077aeef4a00253dedef7003ae73bbd003fffffff"),
                (x"ffffffffff05c0e4a48005ee9edef70009deb817003fffffff"),
                (x"fffffffffff801dbdc9005ef74def7040894f400ffffffffff"),
                (x"fffffffffff801dbdc9005ef74def7040894f400ffffffffff"),
                (x"ffffffffffffc0cbdc9085ef7bdef784097bb01fffffffffff"),
                (x"fffffffffffffe04a6f7bdef7bdef7bdee9483ffffffffffff"),
                (x"fffffffffff79fe63137bdef7bdef7bdd2c679fef7bfffffff"),
                (x"ffffffffde28425f798c4a537bdd294b19ef1421297dffffff"),
                (x"ffffffffde28425f798c4a537bdd294b19ef1421297dffffff"),
                (x"fffffff8a508421f7bdef318c6318cf7bdef0421084befffff"),
                (x"fffffff8a529425f78be2d294652942f8bef1425294befffff"),
                (x"ffffff14210f8bef78be094a3b0ca50f8bef78be08425f7fff"),
                (x"ffffff042179180f782508434650210943ef01847bc21f7fff"),
                (x"ffffff042179180f782508434650210943ef01847bc21f7fff"),
                (x"fffff29421232e9f78212842cb30212843ef26ec210252ffff"),
                (x"ffffff14a5226e929421094a5614a5084252a6e9210a5f7fff"),
                (x"fffffffbde7b2e9294210842129421084252a6ec7bfdefffff"),
                (x"ffffffffff000002942108421f04210842528000003fffffff"),
                (x"ffffffffff000002942108421f04210842528000003fffffff"),
                (x"fffffffffffffff0000708421004842140007fffffffffffff"),
                (x"fffffffffffffff0004210842008421084007fffffffffffff"),
                (x"fffffffffffffff0004238842008423884007fffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc1425280f82942501ffffffffffffffff"),

                -- 1_character_0_3
                (x"fffffffffffffbd739ceef7bdef7bdefffffffffffffffffff"),
                (x"fffffffdce73aa8422ae739d5ad6b573bbdeffffffffffffff"),
                (x"fffffff5ceaa1084210ead6a8bdef7456ae777bfffffffffff"),
                (x"fffffff5ceaa1084210ead6a8bdef7456ae777bfffffffffff"),
                (x"ffffffffbdeb9d5ad6b5ad6b5ad508422b5ab9ddffffffffff"),
                (x"ffffffffffebab5ad5ce756a8bdeb5ad6ae777bfffffffffff"),
                (x"ffffffffbd7550873ab5ab9ceaa108456b5ab9ddffffffffff"),
                (x"ffffffffbd7550873ab5ab9ceaa108456b5ab9ddffffffffff"),
                (x"fffffff5ce75ef5ef6a8ad6ae756b5422b5ad5ddffffffffff"),
                (x"fffffeb9ceaa10eef5d7456ae739cead5d5ad6aeef7fffffff"),
                (x"ffffffffbdaa2bd633ae42115ebbbd756ae73ab573bbffffff"),
                (x"ffffffffbd755dd4a7bd756a8eb9ceebab5af5ddef7fffffff"),
                (x"ffffffffffed7ac4a58ceb9d5af5ce775ce757bdffffffffff"),
                (x"ffffffffffed7ac4a58ceb9d5af5ce775ce757bdffffffffff"),
                (x"ffffffffffebba9bdc002b9ceabbbd777bdeb9ddffffffffff"),
                (x"ffffffffffff537bdc002253d73bbdef7bdef7bdffffffffff"),
                (x"fffffffffff82f7bdc1025ef74f7bd4d3bdef7bdffffffffff"),
                (x"fffffffffff82f7bde1025ef7ba694a77bdef7bfffffffffff"),
                (x"fffffffffff82f7bde1025ef7ba694a77bdef7bfffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694ef7bdef7bfffffffffff"),
                (x"fffffffffff8137bdef7bdef7bb294ef41fff7ffffffffffff"),
                (x"ffffffffffffc09bdef7bdef765294ed3fffffffffffffffff"),
                (x"fffffffffffffe00018c6318cf3def7fbfffffffffffffffff"),
                (x"fffffffffffffe00018c6318cf3def7fbfffffffffffffffff"),
                (x"fffffffffffffffffe94a7bc529421097dffffffffffffffff"),
                (x"ffffffffffffffff7ac3a14a128421087dffffffffffffffff"),
                (x"fffffffffffffff63183294bef14a5084bef7fffffffffffff"),
                (x"fffffffffffffffb5a942fbc4f04212843ef7fffffffffffff"),
                (x"fffffffffffffffb5a942fbc4f04212843ef7fffffffffffff"),
                (x"fffffffffffffffb588565ee9214210843ef7fffffffffffff"),
                (x"fffffffffffffff631e165ee91f821084a007fffffffffffff"),
                (x"ffffffffffffffff78a10252c7f8a52941ffffffffffffffff"),
                (x"ffffffffffffffff78a1094a0f7bde003dffffffffffffffff"),
                (x"ffffffffffffffff78a1094a0f7bde003dffffffffffffffff"),
                (x"ffffffffffffffffffc508421294a52fbdffffffffffffffff"),
                (x"ffffffffffffffffffe2108421084210bfffffffffffffffff"),
                (x"ffffffffffffffffffff01ce739c4207ffffffffffffffffff"),
                (x"ffffffffffffffffffff0084738800ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0084738800ffffffffffffffffffff"),
                (x"ffffffffffffffffffff05284a5000ffffffffffffffffffff"),

                -- 1_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffef7ae739ddeb9ce73bbdeffffffffffffff"),
                (x"fffffffffffffbd73ab5ab9ce756b5ad6ae73bbdffffffffff"),
                (x"fffffffffffffbd73ab5ab9ce756b5ad6ae73bbdffffffffff"),
                (x"ffffffffffff5d5ad517456aead6b5422e8456aeef7fffffff"),
                (x"fffffffffffffae73aa84210eab9ceaa115abbbdffffffffff"),
                (x"ffffffffffff5d5bdd15ab9ce756b575517ba2aeef7fffffff"),
                (x"ffffffffffff5d5bdd15ab9ce756b575517ba2aeef7fffffff"),
                (x"ffffffffbdebaa8ad6b5ad6b5722b5ab915ad6b573bbffffff"),
                (x"fffffff5cead6b5739d5456b572108abaa843ab5ad5ddfffff"),
                (x"ffffffffbd756ae73ab7456ae75ef7ab9d5aa1ddef7bffffff"),
                (x"ffffffffffebab573aa8ad6b5ad508755ce756ae73bfffffff"),
                (x"ffffffffbd756aead6b5aa115756b5756ae73ab573bbffffff"),
                (x"ffffffffbd756aead6b5aa115756b5756ae73ab573bbffffff"),
                (x"fffffff5ceabbaead6aeaa115755ce73aae739ce739dffffff"),
                (x"fffffef7bdef5cead5dd456aeeb9ceef5ce777bd73bbdfffff"),
                (x"ffffffffff076ae73bae456bdebbbd777ae73bbd003fffffff"),
                (x"ffffffffff076aeef7aeab9dd777bd73bae7381d003fffffff"),
                (x"ffffffffff076aeef7aeab9dd777bd73bae7381d003fffffff"),
                (x"fffffffffff81dd73abd777aeaf5ceabbae77400ffffffffff"),
                (x"ffffffffffffc1d73abdeb9ceabab5ab9ddef41fffffffffff"),
                (x"fffffffffffffe0ef5ddeb9d5739ceabbbde83ffffffffffff"),
                (x"fffffffffffffc5003aeef7aeef5ce73ba007bffffffffffff"),
                (x"fffffffffffffc5003aeef7aeef5ce73ba007bffffffffffff"),
                (x"ffffffffffff8a108400ef7bd077bd70001097dfffffffffff"),
                (x"fffffffffff142129425000000000001421087dfffffffffff"),
                (x"fffffffffff14a5f7821294a5294a5284a1084beffffffffff"),
                (x"ffffffffff294bef78210842108421094a108425f7bfffffff"),
                (x"ffffffffff294bef78210842108421094a108425f7bfffffff"),
                (x"ffffffffff014bef78210842108421097c108425f7bfffffff"),
                (x"fffffffffff8000294210842128421097c528425f7bfffffff"),
                (x"fffffffffffffe02942108421f1421084bef14a0ffffffffff"),
                (x"fffffffffffffe02942108421f1421084bef001fffffffffff"),
                (x"fffffffffffffe02942108421f1421084bef001fffffffffff"),
                (x"fffffffffffffe0f78a52fbdef78a5297c007fffffffffffff"),
                (x"fffffffffffffffffc0211ce710842103fffffffffffffffff"),
                (x"ffffffffffffffffffe03c2103800007ffffffffffffffffff"),
                (x"ffffffffffffffffffff05294a03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff05294a03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff0528f183ffffffffffffffffffffff"),

                -- 1_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffdef7bdef7bd739ddef7ffffffffffff"),
                (x"ffffffffffffffdef5cead6b5ab9ce75508455ce73bfffffff"),
                (x"ffffffffffffffdef5cead6b5ab9ce75508455ce73bfffffff"),
                (x"ffffffffffff7aead6a8bdef7456b5721084211573bbffffff"),
                (x"ffffffffffeb9d5ad508456b5ad6b5ad6b5ab9ddef7fffffff"),
                (x"ffffffffffff7aead6b5adef7455ce73ab5ad5ddffffffffff"),
                (x"ffffffffffff7aead6b5adef7455ce73ab5ad5ddffffffffff"),
                (x"ffffffffffeb9d5ad6a84211573ab5ad5c8422aeef7fffffff"),
                (x"ffffffffffebab5ad508ad6ae756b5457b5adeee73bbffffff"),
                (x"ffffffffbd756b573ab5739ce75508bbbae72115739ddfffff"),
                (x"fffffff5cead5cead6aeeb9ddaa1087759ded515ef7fffffff"),
                (x"ffffffffbdebbb5ad5dd739dd455ceef53debaaeef7fffffff"),
                (x"ffffffffbdebbb5ad5dd739dd455ceef53debaaeef7fffffff"),
                (x"ffffffffffef6ae73bae777b5abbbd6312c676bdffffffffff"),
                (x"ffffffffffeb9ddef7aeeb9d5738a5002e94f5ddffffffffff"),
                (x"ffffffffffef7bdef7bdeb9ceea484002f7ba7bfffffffffff"),
                (x"ffffffffffef7bdef689ef7a9bdc84802f7bdc1fffffffffff"),
                (x"ffffffffffef7bdef689ef7a9bdc84802f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7b4a2537bdc84842f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7bda2537bdef7bdef7bdc1fffffffffff"),
                (x"fffffffffffffbf003bda3197bdef7bdef7ba41fffffffffff"),
                (x"fffffffffffffffffe9da528cbdef7bdee9483ffffffffffff"),
                (x"fffffffffffffffffe9da528cbdef7bdee9483ffffffffffff"),
                (x"ffffffffffffffffffde294a26318c6300007fffffffffffff"),
                (x"ffffffffffffffffffc508425f7bde103fffffffffffffffff"),
                (x"fffffffffffffff000a10842529421a101ffffffffffffffff"),
                (x"fffffffffffffff000a1084251fbde10d9ffffffffffffffff"),
                (x"fffffffffffffff000a1084251fbde10d9ffffffffffffffff"),
                (x"fffffffffffffe0f78a1094a123129b859ffffffffffffffff"),
                (x"fffffffffffffe0297c508421232f7b819ffffffffffffffff"),
                (x"ffffffffffffffe297c5294a11b129b805ffffffffffffffff"),
                (x"fffffffffffffe5294bef14a528d8c0085ffffffffffffffff"),
                (x"fffffffffffffe5294bef14a528d8c0085ffffffffffffffff"),
                (x"ffffffffffffffef78a5f7bdef00001081ffffffffffffffff"),
                (x"ffffffffffffffef7800f14a52fbde103fffffffffffffffff"),
                (x"fffffffffffffe0108f0388420004210bfffffffffffffffff"),
                (x"fffffffffffffff000f081ce0f8294a53fffffffffffffffff"),
                (x"fffffffffffffff000f081ce0f8294a53fffffffffffffffff"),
                (x"fffffffffffffffa5294a1080fffffffffffffffffffffffff"),

                -- 1_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffef7ae739ceef5ce73bbdeffffffffffffff"),
                (x"ffffffffffff7ae73ab5ad6b5739cead6ae777bfffffffffff"),
                (x"ffffffffffff7ae73ab5ad6b5739cead6ae777bfffffffffff"),
                (x"ffffffffffebab5422e8456b5abab545d15ad5ddffffffffff"),
                (x"ffffffffffff7aead508ab9ceab908422ae73bbfffffffffff"),
                (x"ffffffffffebaa8bdd15756b5777bd75517bd5ddffffffffff"),
                (x"ffffffffffebaa8bdd15756b5777bd75517bd5ddffffffffff"),
                (x"ffffffffbd756b5ad50ead6a8775ceabab5aa2aeef7bffffff"),
                (x"fffffff5cead6ae422ae42108777bd455ce756b5ad5ddfffff"),
                (x"ffffffffbdef5c8ad6ae45ef7777bd45dce73ab573bbffffff"),
                (x"ffffffffff73ab573aaeaa115733bd722bdeb9d5ef7fffffff"),
                (x"ffffffffbd756aead6ae756b57258ced6ae775ce73bbffffff"),
                (x"ffffffffbd756aead6ae756b57258ced6ae775ce73bbffffff"),
                (x"fffffffdceab9cead5ddeb9d5edd29ebaae775ce739ddfffff"),
                (x"fffffff7bd777ae73bac677aeedef7675d5af5ddef7bdeffff"),
                (x"ffffffffff077aeef4a00253dedef7003ae73bbd003fffffff"),
                (x"ffffffffff05c0e4a48005ee9edef70009deb817003fffffff"),
                (x"ffffffffff05c0e4a48005ee9edef70009deb817003fffffff"),
                (x"fffffffffff801dbdc9005ef74def7040894f400ffffffffff"),
                (x"ffffffffffffc0cbdc9085ef7bdef784097bb01fffffffffff"),
                (x"fffffffffffffe04a6f7bdef7bdef7bdee9483ffffffffffff"),
                (x"ffffffffffff8be63137bdef7bdef7bdd2c678beffffffffff"),
                (x"ffffffffffff8be63137bdef7bdef7bdd2c678beffffffffff"),
                (x"ffffffffff28425f798c4a537bdd294b18528425f7bfffffff"),
                (x"ffffffffde28421294bef318c6318cf7bc108421297dffffff"),
                (x"fffffff8a529425f78252d29465294294a1094a1297dffffff"),
                (x"fffffff8a5294be294a1094a3b0ca5097c528425297dffffff"),
                (x"fffffff8a5294be294a1094a3b0ca5097c528425297dffffff"),
                (x"ffffff94a5297c0294a5094b4650a50846420421297dffffff"),
                (x"fffffff88420c0008421294acb30a52b2e9490a1f7bfffffff"),
                (x"ffffffbc634bc1e0842108421614210b2f7b8ca5003fffffff"),
                (x"ffffff818c4b3fe2942108421294210952948ca0ffffffffff"),
                (x"ffffff818c4b3fe2942108421294210952948ca0ffffffffff"),
                (x"fffffffc00003fff78a52fbde078a52fbc00001fffffffffff"),
                (x"fffffffffffffff0000211ce7388421084007fffffffffffff"),
                (x"fffffffffffffffffc023c210388421001ffffffffffffffff"),
                (x"ffffffffffffffffffe081ce21000007ffffffffffffffffff"),
                (x"ffffffffffffffffffe081ce21000007ffffffffffffffffff"),
                (x"ffffffffffffffffffff05294203ffffffffffffffffffffff"),

                -- 1_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffbd739ceef7bdef7bdefffffffffffffffffff"),
                (x"fffffffdce73aa8422ae739d5ad6b573bbdeffffffffffffff"),
                (x"fffffffdce73aa8422ae739d5ad6b573bbdeffffffffffffff"),
                (x"fffffff5ceaa1084210ead6a8bdef7456ae777bfffffffffff"),
                (x"ffffffffbdeb9d5ad6b5ad6b5ad508422b5ab9ddffffffffff"),
                (x"ffffffffffebab5ad5ce756a8bdeb5ad6ae777bfffffffffff"),
                (x"ffffffffffebab5ad5ce756a8bdeb5ad6ae777bfffffffffff"),
                (x"ffffffffbd7550873ab5ab9ceaa108456b5ab9ddffffffffff"),
                (x"fffffff5ce75ef5ef6a8ad6ae756b5422b5ad5ddffffffffff"),
                (x"fffffeb9ceaa10eef5d7456ae739cead5d5ad6aeef7fffffff"),
                (x"ffffffffbdaa2bd633ae42115ebbbd756ae73ab573bbffffff"),
                (x"ffffffffbd755dd4a7bd756a8eb9ceebab5af5ddef7fffffff"),
                (x"ffffffffbd755dd4a7bd756a8eb9ceebab5af5ddef7fffffff"),
                (x"ffffffffffed7ac4a58ceb9d5af5ce775ce757bdffffffffff"),
                (x"ffffffffffebba9bdc002b9ceabbbd777bdeb9ddffffffffff"),
                (x"ffffffffffff537bdc002253d73bbdef7bdef7bdffffffffff"),
                (x"fffffffffff82f7bdc1025ef74f7bd4d3bdef7bdffffffffff"),
                (x"fffffffffff82f7bdc1025ef74f7bd4d3bdef7bdffffffffff"),
                (x"fffffffffff82f7bde1025ef7ba694a77bdef7bfffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694ef7bdef7bfffffffffff"),
                (x"fffffffffff8137bdef7bdef7bb294ef41fff7ffffffffffff"),
                (x"ffffffffffffc09bdef7bdef765294ed3fffffffffffffffff"),
                (x"ffffffffffffc09bdef7bdef765294ed3fffffffffffffffff"),
                (x"fffffffffffffe00018c6318cf14a510bfffffffffffffffff"),
                (x"fffffffffffffffffc1ef7bde284212fbfffffffffffffffff"),
                (x"fffffffffffffff00094094a5284210941ffffffffffffffff"),
                (x"fffffffffffffff6307ef7bc3284210941ffffffffffffffff"),
                (x"fffffffffffffff6307ef7bc3284210941ffffffffffffffff"),
                (x"fffffffffffffff630374b18409421097c007fffffffffffff"),
                (x"fffffffffffffff63017bb184084212f8a007fffffffffffff"),
                (x"ffffffffffffffff78174b183094a52f8bef7fffffffffffff"),
                (x"ffffffffffffffff7bc060c65297def14a52ffffffffffffff"),
                (x"ffffffffffffffff7bc060c65297def14a52ffffffffffffff"),
                (x"fffffffffffffff003de0001ef7bde297def7fffffffffffff"),
                (x"fffffffffffffffffc02f7bc5297de003def7fffffffffffff"),
                (x"fffffffffffffffffc4210000108e781c4007fffffffffffff"),
                (x"fffffffffffffffffe94a001f01e1081c1ffffffffffffffff"),
                (x"fffffffffffffffffe94a001f01e1081c1ffffffffffffffff"),
                (x"fffffffffffffffffffffffff01294a501ffffffffffffffff"),

                -- 1_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffef7ae739ddeb9ce73bbdeffffffffffffff"),
                (x"fffffffffffffbd73ab5ab9ce756b5ad6ae73bbdffffffffff"),
                (x"fffffffffffffbd73ab5ab9ce756b5ad6ae73bbdffffffffff"),
                (x"ffffffffffff5d5ad517456aead6b5422e8456aeef7fffffff"),
                (x"fffffffffffffae73aa84210eab9ceaa115abbbdffffffffff"),
                (x"ffffffffffff5d5bdd15ab9ce756b575517ba2aeef7fffffff"),
                (x"ffffffffffff5d5bdd15ab9ce756b575517ba2aeef7fffffff"),
                (x"ffffffffbdebaa8ad6b5ad6b5722b5ab915ad6b573bbffffff"),
                (x"fffffff5cead6b5739d5456b572108abaa843ab5ad5ddfffff"),
                (x"ffffffffbd756ae73ab7456ae75ef7ab9d5aa1ddef7bffffff"),
                (x"ffffffffffebab573aa8ad6b5ad508755ce756ae73bfffffff"),
                (x"ffffffffbd756aead6b5aa115756b5756ae73ab573bbffffff"),
                (x"ffffffffbd756aead6b5aa115756b5756ae73ab573bbffffff"),
                (x"fffffff5ceabbaead6aeaa115755ce73aae739ce739dffffff"),
                (x"fffffef7bdef5cead5dd456aeeb9ceef5ce777bd73bbdfffff"),
                (x"ffffffffff076ae73bae456bdebbbd777ae73bbd003fffffff"),
                (x"ffffffffff076aeef7aeab9dd777bd73bae7381d003fffffff"),
                (x"ffffffffff076aeef7aeab9dd777bd73bae7381d003fffffff"),
                (x"fffffffffff81dd73abd777aeaf5ceabbae77400ffffffffff"),
                (x"ffffffffffffc1d73abdeb9ceabab5ab9ddef41fffffffffff"),
                (x"fffffffffffffe0ef5ddeb9d5739ceabbbde83ffffffffffff"),
                (x"fffffffffffffe2003aeef7aeef5ce73ba0017dfffffffffff"),
                (x"fffffffffffffe2003aeef7aeef5ce73ba0017dfffffffffff"),
                (x"fffffffffffffc508400ef7bd077bd70001084beffffffffff"),
                (x"fffffffffffffc10842500000000000142528425f7bfffffff"),
                (x"ffffffffffff8a1084a1294a5294a52843ef14a5f7bfffffff"),
                (x"fffffffffff1421084a508421084210843ef78a5297fffffff"),
                (x"fffffffffff1421084a508421084210843ef78a5297fffffff"),
                (x"fffffffffff1421087c508421084210843ef78a5003fffffff"),
                (x"fffffffffff1421297c508421284210842528000ffffffffff"),
                (x"fffffffffff80a5f78a108425f042108425283ffffffffffff"),
                (x"ffffffffffffc00f78a108425f042108425283ffffffffffff"),
                (x"ffffffffffffc00f78a108425f042108425283ffffffffffff"),
                (x"fffffffffffffff003c5294bef7bde294a2103ffffffffffff"),
                (x"ffffffffffffffffffe01084211ce71081ffffffffffffffff"),
                (x"ffffffffffffffffffff000003c210383fffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a529407ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a529407ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe01be9407ffffffffffffffffff"),

                -- 1_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffdef7bdef7bd739ddef7ffffffffffff"),
                (x"ffffffffffffffdef5cead6b5ab9ce75508455ce73bfffffff"),
                (x"ffffffffffffffdef5cead6b5ab9ce75508455ce73bfffffff"),
                (x"ffffffffffff7aead6a8bdef7456b5721084211573bbffffff"),
                (x"ffffffffffeb9d5ad508456b5ad6b5ad6b5ab9ddef7fffffff"),
                (x"ffffffffffff7aead6b5adef7455ce73ab5ad5ddffffffffff"),
                (x"ffffffffffff7aead6b5adef7455ce73ab5ad5ddffffffffff"),
                (x"ffffffffffeb9d5ad6a84211573ab5ad5c8422aeef7fffffff"),
                (x"ffffffffffebab5ad508ad6ae756b5457b5adeee73bbffffff"),
                (x"ffffffffbd756b573ab5739ce75508bbbae72115739ddfffff"),
                (x"fffffff5cead5cead6aeeb9ddaa1087759ded515ef7fffffff"),
                (x"ffffffffbdebbb5ad5dd739dd455ceef53debaaeef7fffffff"),
                (x"ffffffffbdebbb5ad5dd739dd455ceef53debaaeef7fffffff"),
                (x"ffffffffffef6ae73bae777b5abbbd6312c676bdffffffffff"),
                (x"ffffffffffeb9ddef7aeeb9d5738a5002e94f5ddffffffffff"),
                (x"ffffffffffef7bdef7bdeb9ceea484002f7ba7bfffffffffff"),
                (x"ffffffffffef7bdef689ef7a9bdc84802f7bdc1fffffffffff"),
                (x"ffffffffffef7bdef689ef7a9bdc84802f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7b4a2537bdc84842f7bdc1fffffffffff"),
                (x"ffffffffffff7bdef7bda2537bdef7bdef7bdc1fffffffffff"),
                (x"fffffffffffffbf003bda3197bdef7bdef7ba41fffffffffff"),
                (x"fffffffffffffffffe9da528cbdef7bdee9483ffffffffffff"),
                (x"fffffffffffffffffe9da528cbdef7bdee9483ffffffffffff"),
                (x"fffffffffffffff003c52fbde6318c6300007fffffffffffff"),
                (x"fffffffffffffe0f78a108425f7a94a53fffffffffffffffff"),
                (x"ffffffffffffffe2942128421f0463b0e9ffffffffffffffff"),
                (x"ffffffffffffc0508425f14a1f06946328c67fffffffffffff"),
                (x"ffffffffffffc0508425f14a1f06946328c67fffffffffffff"),
                (x"ffffffffffffc05084a10fbc5284a5a5bc94b3ffffffffffff"),
                (x"ffffffffffffc052942109083f1421233c9483ffffffffffff"),
                (x"fffffffffffffe0294a120c77678a5a17c007fffffffffffff"),
                (x"fffffffffffffe0f78a52319767821097dffffffffffffffff"),
                (x"fffffffffffffe0f78a52319767821097dffffffffffffffff"),
                (x"fffffffffffffe2000021b189014212fbdffffffffffffffff"),
                (x"fffffffffffffe210842100021084210bfffffffffffffffff"),
                (x"fffffffffffffff108400000011ce738bfffffffffffffffff"),
                (x"fffffffffffffff00294a7fe01084213c1ffffffffffffffff"),
                (x"fffffffffffffff00294a7fe01084213c1ffffffffffffffff"),
                (x"fffffffffffffffffffffffffa5294a101ffffffffffffffff"),

                -- 1_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffef7ae739ceef5ce73bbdeffffffffffffff"),
                (x"ffffffffffff7ae73ab5ad6b5739cead6ae777bfffffffffff"),
                (x"ffffffffffff7ae73ab5ad6b5739cead6ae777bfffffffffff"),
                (x"ffffffffffebab5422e8456b5abab545d15ad5ddffffffffff"),
                (x"ffffffffffff7aead508ab9ceab908422ae73bbfffffffffff"),
                (x"ffffffffffebaa8bdd15756b5777bd75517bd5ddffffffffff"),
                (x"ffffffffffebaa8bdd15756b5777bd75517bd5ddffffffffff"),
                (x"ffffffffbd756b5ad50ead6a8775ceabab5aa2aeef7bffffff"),
                (x"fffffff5cead6ae422ae42108777bd455ce756b5ad5ddfffff"),
                (x"ffffffffbdef5c8ad6ae45ef7777bd45dce73ab573bbffffff"),
                (x"ffffffffff73ab573aaeaa115733bd722bdeb9d5ef7fffffff"),
                (x"ffffffffbd756aead6ae756b57258ced6ae775ce73bbffffff"),
                (x"ffffffffbd756aead6ae756b57258ced6ae775ce73bbffffff"),
                (x"fffffffdceab9cead5ddeb9d5edd29ebaae775ce739ddfffff"),
                (x"fffffff7bd777ae73bac677aeedef7675d5af5ddef7bdeffff"),
                (x"ffffffffff077aeef4a00253dedef7003ae73bbd003fffffff"),
                (x"ffffffffff05c0e4a48005ee9edef70009deb817003fffffff"),
                (x"ffffffffff05c0e4a48005ee9edef70009deb817003fffffff"),
                (x"fffffffffff801dbdc9005ef74def7040894f400ffffffffff"),
                (x"ffffffffffffc0cbdc9085ef7bdef784097bb01fffffffffff"),
                (x"fffffffffffffe04a6f7bdef7bdef7bdee9483ffffffffffff"),
                (x"ffffffffffff8be63137bdef7bdef7bdd2c678beffffffffff"),
                (x"ffffffffffff8be63137bdef7bdef7bdd2c678beffffffffff"),
                (x"fffffffffff14212958c4a537bdd294b19ef1421297fffffff"),
                (x"ffffffffde28421087def318c6318cf78a528421297dffffff"),
                (x"ffffffffde284a5084a52d294652942943ef1425294befffff"),
                (x"ffffffffde29421297c5094a3b0ca5084a52f8a5294befffff"),
                (x"ffffffffde29421297c5094a3b0ca5084a52f8a5294befffff"),
                (x"ffffffffde2842121061094b4650a5094a5283c5294a5fffff"),
                (x"fffffffffff04a44a6ec294acb30a528421080032109efffff"),
                (x"ffffffffff014a3bdeec0842560421084210f80f4a46ffffff"),
                (x"fffffffffff80a34a5250842528421084252fbec4a580fffff"),
                (x"fffffffffff80a34a5250842528421084252fbec4a580fffff"),
                (x"ffffffffffffc00003de294be07bde294bef7fe00001ffffff"),
                (x"fffffffffffffff000421084239ce71080007fffffffffffff"),
                (x"fffffffffffffffffc00108423c2103881ffffffffffffffff"),
                (x"ffffffffffffffffffff00000108e7803fffffffffffffffff"),
                (x"ffffffffffffffffffff00000108e7803fffffffffffffffff"),
                (x"ffffffffffffffffffffffff42529407ffffffffffffffffff"),

                -- 1_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffbd739ceef7bdef7bdefffffffffffffffffff"),
                (x"fffffffdce73aa8422ae739d5ad6b573bbdeffffffffffffff"),
                (x"fffffffdce73aa8422ae739d5ad6b573bbdeffffffffffffff"),
                (x"fffffff5ceaa1084210ead6a8bdef7456ae777bfffffffffff"),
                (x"ffffffffbdeb9d5ad6b5ad6b5ad508422b5ab9ddffffffffff"),
                (x"ffffffffffebab5ad5ce756a8bdeb5ad6ae777bfffffffffff"),
                (x"ffffffffffebab5ad5ce756a8bdeb5ad6ae777bfffffffffff"),
                (x"ffffffffbd7550873ab5ab9ceaa108456b5ab9ddffffffffff"),
                (x"fffffff5ce75ef5ef6a8ad6ae756b5422b5ad5ddffffffffff"),
                (x"fffffeb9ceaa10eef5d7456ae739cead5d5ad6aeef7fffffff"),
                (x"ffffffffbdaa2bd633ae42115ebbbd756ae73ab573bbffffff"),
                (x"ffffffffbd755dd4a7bd756a8eb9ceebab5af5ddef7fffffff"),
                (x"ffffffffbd755dd4a7bd756a8eb9ceebab5af5ddef7fffffff"),
                (x"ffffffffffed7ac4a58ceb9d5af5ce775ce757bdffffffffff"),
                (x"ffffffffffebba9bdc002b9ceabbbd777bdeb9ddffffffffff"),
                (x"ffffffffffff537bdc002253d73bbdef7bdef7bdffffffffff"),
                (x"fffffffffff82f7bdc1025ef74f7bd4d3bdef7bdffffffffff"),
                (x"fffffffffff82f7bdc1025ef74f7bd4d3bdef7bdffffffffff"),
                (x"fffffffffff82f7bde1025ef7ba694a77bdef7bfffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694ef7bdef7bfffffffffff"),
                (x"fffffffffff8137bdef7bdef7bb294ef41fff7ffffffffffff"),
                (x"ffffffffffffc09bdef7bdef765294ed3fffffffffffffffff"),
                (x"ffffffffffffc09bdef7bdef765294ed3fffffffffffffffff"),
                (x"fffffffffffffe00018c6318cf78e73f81ffffffffffffffff"),
                (x"fffffffffffffffffe94a7bde28421097c007fffffffffffff"),
                (x"fffffffffffffffa50761843e084a5084bef7fffffffffffff"),
                (x"fffffffffffffeca518ca043e097de28425283ffffffffffff"),
                (x"fffffffffffffeca518ca043e097de28425283ffffffffffff"),
                (x"ffffffffffffd89f7ad4284252f82109425283ffffffffffff"),
                (x"ffffffffffffc09f7984094be19021084a5283ffffffffffff"),
                (x"fffffffffffffe0f78af2fbccb8c84094a007fffffffffffff"),
                (x"ffffffffffffffff78a10fbccbb084297c007fffffffffffff"),
                (x"ffffffffffffffff78a10fbccbb084297c007fffffffffffff"),
                (x"ffffffffffffffff7bc5094a04b063f000217fffffffffffff"),
                (x"fffffffffffffffffc4210842100421084217fffffffffffff"),
                (x"fffffffffffffffffc4739ce2000000085ffffffffffffffff"),
                (x"fffffffffffffff001e21084207e94a501ffffffffffffffff"),
                (x"fffffffffffffff001e21084207e94a501ffffffffffffffff"),
                (x"fffffffffffffff00094a5280fffffffffffffffffffffffff"),

                -- 2_character_0_0
                (x"ffffffffffffffffffee739ce739ce73bfffffffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5756ae77fffffffffffff"),
                (x"ffffffffffffdd5ad517ad6a8aa2b5aa115ad5dfffffffffff"),
                (x"ffffffffffffdd5ad517ad6a8aa2b5aa115ad5dfffffffffff"),
                (x"fffffffffffbaa8422a8bd6b7422b5422b5aa2aeffffffffff"),
                (x"fffffffffffd51742115ba117455084550842115ffffffffff"),
                (x"ffffffffff722f742108421084550842108422f573bfffffff"),
                (x"ffffffffff722f742108421084550842108422f573bfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d1573bfffffff"),
                (x"ffffffffbdadee8422f7ba117ba2f7bdef7ba115ad7bffffff"),
                (x"ffffffffbd45d0842108bdef7bdef7bdd0842115ad7bffffff"),
                (x"fffffffdce42108421084211742108ba2a8422a8ad5dffffff"),
                (x"fffffff6b542108421084210842108422a8422a8ad6bdfffff"),
                (x"fffffff6b542108421084210842108422a8422a8ad6bdfffff"),
                (x"fffffff50845508422a84210842108422a8422a873abdfffff"),
                (x"ffffffb90845508422a84210842108422a8422a873aaefffff"),
                (x"ffffffb90845515422a8456a8aa108422a84551573aaefffff"),
                (x"fffffff6b543915422b5456a8aa108455c84551573abdfffff"),
                (x"fffffff6b543915422b5456a8aa108455c84551573abdfffff"),
                (x"fffffff5ce43ab5422b5456a8aa108455c84390ead5ddfffff"),
                (x"ffffffffbdaf6ae422ae456a8ad508abab5abaaead7bffffff"),
                (x"ffffffffff077aead6aeab9d5756b5776ae73bbd003fffffff"),
                (x"ffffffffffffe9def5cc777aeebbbdeb3bdef69fffffffffff"),
                (x"ffffffffffffe9def5cc777aeebbbdeb3bdef69fffffffffff"),
                (x"fffffffffffd0a5631c42318c6318c211cc61194ffffffffff"),
                (x"ffffffffffa1484a5084210842108421094a1085a53fffffff"),
                (x"ffffffffff71485a50a42042108421210b4a148573bfffffff"),
                (x"fffffffe94094a500284210842108421280014a50869ffffff"),
                (x"fffffffe94094a500284210842108421280014a50869ffffff"),
                (x"ffffffd1ce2848e0028521084210842168003881295d4fffff"),
                (x"ffffffd084094a0ffca42042108421210bff80a508494fffff"),
                (x"fffffffc007048000084204210842121080000817381ffffff"),
                (x"fffffffc004a41fa51c42042108421211d4a7c094a41ffffff"),
                (x"fffffffc004a41fa51c42042108421211d4a7c094a41ffffff"),
                (x"ffffffffff003ffa53bef7bdef7bdef7bb4a7fe0003fffffff"),
                (x"fffffffffffffffa53bdf7bdef7bdef77b4a7fffffffffffff"),
                (x"fffffffffffffff0019df77ac033bdf758007fffffffffffff"),
                (x"fffffffffffffffffc1d1f7a0f83bd1f41ffffffffffffffff"),
                (x"fffffffffffffffffc1d1f7a0f83bd1f41ffffffffffffffff"),
                (x"fffffffffffffffffc0cb3180f818cb301ffffffffffffffff"),

                -- 2_character_0_1
                (x"fffffffffffffffffdce739d5ad6b5739dffffffffffffffff"),
                (x"fffffffffffffee73aa845ef7ba2b5aa2ae73bffffffffffff"),
                (x"ffffffffffffdd542117bdef7bdef7ba10845ebfffffffffff"),
                (x"ffffffffffffdd542117bdef7bdef7ba10845ebfffffffffff"),
                (x"fffffffffffbaa8ad508456b5ad508bdd15aa2eeffffffffff"),
                (x"ffffffffff7551542115aa108ba2b5aa2e8456f5ffffffffff"),
                (x"ffffffffff756a8422a842117455294bab5ad5d573bfffffff"),
                (x"ffffffffff756a8422a842117455294bab5ad5d573bfffffff"),
                (x"fffffffdcead6a8ad508aa108aa6f7bdd2e7393573bfffffff"),
                (x"fffffffdcead50842115adee8adef7bdef7bdd3573bfffffff"),
                (x"fffffffdcead5154211545ef54def7bdef7bdd2effffffffff"),
                (x"ffffffbab5ab915422b545ef5bdef7bdef7bdd9dffffffffff"),
                (x"ffffffbab5ab90e422ae42115ba58c632f7bdc1fffffffffff"),
                (x"ffffffbab5ab90e422ae42115ba58c632f7bdc1fffffffffff"),
                (x"ffffffbab57550e422aeaa115ba4a5002f7bdc1fffffffffff"),
                (x"fffffff6b5756aead5d7aa10eba484002f7bdc1fffffffffff"),
                (x"fffffff6b5756aead7a97210ebdc8439ef7bdc1fffffffffff"),
                (x"fffffff5ceebaaead7b4756aebdc8491ef7bdc1fffffffffff"),
                (x"fffffff5ceebaaead7b4756aebdc8491ef7bdc1fffffffffff"),
                (x"ffffffffbda75cead7bd739c9bdef7bdef7bdc1fffffffffff"),
                (x"fffffffffffd3ae73bbda39c9bdef7bdef7ba41fffffffffff"),
                (x"ffffffffffffff4ef694a528c4def7bdee9483ffffffffffff"),
                (x"fffffffffffffffffe942d28e6318c6300007fffffffffffff"),
                (x"fffffffffffffffffe942d28e6318c6300007fffffffffffff"),
                (x"fffffffffffffffffe8409084a1694a1294a13ffffffffffff"),
                (x"fffffffffffffffa50a409094210a50ba9ef53ffffffffffff"),
                (x"fffffffffffffffa50a421094a042123a9ef53ffffffffffff"),
                (x"fffffffffffffffa50a4214b4290210929ef7fffffffffffff"),
                (x"fffffffffffffffa50a4214b4290210929ef7fffffffffffff"),
                (x"ffffffffffffff473a8529094290842929ef53ffffffffffff"),
                (x"ffffffffffffff42948109085290212869ef53ffffffffffff"),
                (x"ffffffffffffff4738a52108520421207bef53ffffffffffff"),
                (x"fffffffffffffffa502120004090840f7bef53ffffffffffff"),
                (x"fffffffffffffffa502120004090840f7bef53ffffffffffff"),
                (x"fffffffffffffffa5189b801de8421f7ba007fffffffffffff"),
                (x"fffffffffffffffffc00077bdefbdeef41ffffffffffffffff"),
                (x"ffffffffffffffffffe00318c63000003fffffffffffffffff"),
                (x"ffffffffffffffffffff0319ef7400ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0319ef7400ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0318cb3000ffffffffffffffffffff"),

                -- 2_character_0_2
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5ad5ce77fffffffffffff"),
                (x"ffffffffffffdd5ad6a8bdef5aa2f7ba115ab9dfffffffffff"),
                (x"ffffffffffffdd5ad6a8bdef5aa2f7ba115ab9dfffffffffff"),
                (x"fffffffffffbaa8bdef74211745ef7bdee8422aeffffffffff"),
                (x"fffffffffffd50842108bdee845ef7456a842115ffffffffff"),
                (x"ffffffffff756a8bdef742117422b5aa2f7ba11573bfffffff"),
                (x"ffffffffff756a8bdef742117422b5aa2f7ba11573bfffffff"),
                (x"ffffffffff756b5ad6a8bb9d545508bdd08456b573bfffffff"),
                (x"ffffffffbdad508ad5c9ba52eab929ba5d5aa2b5ad7bffffff"),
                (x"ffffffffbdaa11773937bdef7bdef7bdd2e72115ad7bffffff"),
                (x"fffffffdce456f573af7bdef7bdef7bdeee7550ead5dffffff"),
                (x"fffffff5ceabaf573af7bdef7bdef7bdeee756eead5ddfffff"),
                (x"fffffff5ceabaf573af7bdef7bdef7bdeee756eead5ddfffff"),
                (x"fffffff5ceaf50e4a58c65ef7bdef7631894bafd73abdfffff"),
                (x"fffffff6b57250ebdca005ef7bdef7000b7bb90973abdfffff"),
                (x"fffffff6b575eaebdc8005ef7bdef700097bbab773abdfffff"),
                (x"fffffff6b5e82bdbdc873def7bdef739c97bf6a0ef5ddfffff"),
                (x"fffffff6b5e82bdbdc873def7bdef739c97bf6a0ef5ddfffff"),
                (x"fffffff5cee81c0bdc923def7bdef73c897b81c0ef5ddfffff"),
                (x"fffffff5cee83a04a6f7bdef7bdef7bdee9483a0ef5ddfffff"),
                (x"ffffffffbd07c0063137bdef7bdef7bdd2c6001f003bffffff"),
                (x"ffffffffffffe85a500c4a537bdd294b014a329fffffffffff"),
                (x"ffffffffffffe85a500c4a537bdd294b014a329fffffffffff"),
                (x"fffffffffffd0a4295c56318c6318c615c5290b4ffffffffff"),
                (x"ffffffffffa1484a50842109ef788421094a1085a53fffffff"),
                (x"ffffffffff71485a50a10843ef7821084b4a148573bfffffff"),
                (x"fffffffe94094a5000a40843ef7821090a0014a50869ffffff"),
                (x"fffffffe94094a5000a40843ef7821090a0014a50869ffffff"),
                (x"ffffffd1ce2848e002852109ef78842168003881295d4fffff"),
                (x"ffffffd084094a0ffca42109ef7884210bff80a508494fffff"),
                (x"fffffffc0070480000840843ef782109080000817381ffffff"),
                (x"fffffffc004a41fa508108434ed02108494a7c094a41ffffff"),
                (x"fffffffc004a41fa508108434ed02108494a7c094a41ffffff"),
                (x"ffffffffff003ffa53a40d29def694093b4a7fe0003fffffff"),
                (x"fffffffffffffffa53bdf7bddef7def77b4a7fffffffffffff"),
                (x"fffffffffffffff0019ef77ac033bdf798007fffffffffffff"),
                (x"fffffffffffffffffc1d1f7a0f83bd1f41ffffffffffffffff"),
                (x"fffffffffffffffffc1d1f7a0f83bd1f41ffffffffffffffff"),
                (x"fffffffffffffffffc0cb3180f818cb301ffffffffffffffff"),

                -- 2_character_0_3
                (x"fffffffffffffff739cead6b5ab9ce73bfffffffffffffffff"),
                (x"ffffffffffffdcead515aa117bdd08455ce77fffffffffffff"),
                (x"fffffffffffd6e842117bdef7bdef7ba115abbffffffffffff"),
                (x"fffffffffffd6e842117bdef7bdef7ba115abbffffffffffff"),
                (x"ffffffffff75d15422f7456b5ad508422a8455dfffffffffff"),
                (x"ffffffffffadea8bdd15aa117422b5aa115aa2aeffffffffff"),
                (x"fffffffdceabab5ad5c94d6a8ba10845508456aeffffffffff"),
                (x"fffffffdceabab5ad5c94d6a8ba10845508456aeffffffffff"),
                (x"fffffffdceaa5ce4a6f7ba535422b5422a8456b573bfffffff"),
                (x"fffffffdceaa6f7bdef7bdef545eb5aa108422b573bfffffff"),
                (x"ffffffffff726f7bdef7bdee9add08aa115aa2b573bfffffff"),
                (x"ffffffffffeb2f7bdef7bdef7add08ad515aa1d5ad5dffffff"),
                (x"fffffffffff82f7bdd8c62537aa1087550e721d5ad5dffffff"),
                (x"fffffffffff82f7bdd8c62537aa1087550e721d5ad5dffffff"),
                (x"fffffffffff82f7bdc002a537aa2b57550e722aead5dffffff"),
                (x"fffffffffff82f7bdc0022537722b5bbaae756aead7bffffff"),
                (x"fffffffffff82f7bdce725ef7721ce4f6ae756aead7bffffff"),
                (x"fffffffffff82f7bdcf225ef7755cea76ae755dd73bbffffff"),
                (x"fffffffffff82f7bdcf225ef7755cea76ae755dd73bbffffff"),
                (x"fffffffffff82f7bdef7bdef74b9ceef6ae73bb4ef7fffffff"),
                (x"fffffffffff8137bdef7bdef74ba94ef5ce7769fffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a53b4a7fffffffffffff"),
                (x"fffffffffffffe00018c6318c7518ca53fffffffffffffffff"),
                (x"fffffffffffffe00018c6318c7518ca53fffffffffffffffff"),
                (x"ffffffffffffc94a5094a14b421021253fffffffffffffffff"),
                (x"ffffffffffffe9ea51c129084a10212169ffffffffffffffff"),
                (x"ffffffffffffe9ea51c408434a10842169ffffffffffffffff"),
                (x"ffffffffffffffea508109085a14842169ffffffffffffffff"),
                (x"ffffffffffffffea508109085a14842169ffffffffffffffff"),
                (x"ffffffffffffe9ea508521085a10a52d1d4a7fffffffffffff"),
                (x"ffffffffffffe9ea50250908529021090b4a7fffffffffffff"),
                (x"ffffffffffffe9eef4240842429084295d4a7fffffffffffff"),
                (x"ffffffffffffe9eef7a121081200840869ffffffffffffffff"),
                (x"ffffffffffffe9eef7a121081200840869ffffffffffffffff"),
                (x"fffffffffffffe0ef7de0843de82f74b29ffffffffffffffff"),
                (x"fffffffffffffff003bdf7bddef400003fffffffffffffffff"),
                (x"fffffffffffffffffc000318c6300007ffffffffffffffffff"),
                (x"ffffffffffffffffffff077bef3000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff077bef3000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff0319663000ffffffffffffffffffff"),

                -- 2_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce73bfffffffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5756ae77fffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5756ae77fffffffffffff"),
                (x"ffffffffffffdd5ad517ad6a8aa2b5aa115ad5dfffffffffff"),
                (x"fffffffffffbaa8422a8bd6b7422b5422b5aa2aeffffffffff"),
                (x"fffffffffffd51742115ba117455084550842115ffffffffff"),
                (x"fffffffffffd51742115ba117455084550842115ffffffffff"),
                (x"ffffffffff722f742108421084550842108422f573bfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d1573bfffffff"),
                (x"ffffffffbdadee8422f7ba117ba2f7bdef7ba115ad7bffffff"),
                (x"ffffffffbd45d0842108bdef7bdef7bdd0842115ad5dffffff"),
                (x"fffffffdce42108421084211742108ba108422a8ad6bdfffff"),
                (x"fffffffdce42108421084211742108ba108422a8ad6bdfffff"),
                (x"fffffff5ce42108421084210842108422a8422a873aaefffff"),
                (x"fffffff6b542108421084210842108422a8422a873ab5fffff"),
                (x"ffffffbab545508421084210842108422a8421c8ad5d577fff"),
                (x"ffffffbab545508421154210845508421d5aa1d5421d5effff"),
                (x"ffffffbab545508421154210845508421d5aa1d5421d5effff"),
                (x"fffffffdce422a8ad5154211545508421d5aa1ce421ceeffff"),
                (x"ffffffffbdaa1c8ad515aa115456b5421ce755cead5ddfffff"),
                (x"ffffffffffed5d5ad51572115455ce455ce755ddef41ffffff"),
                (x"ffffffffffff7bd73ab5756aead7bdabbae73bbfffffffffff"),
                (x"ffffffffffff7bd73ab5756aead7bdabbae73bbfffffffffff"),
                (x"ffffffffffffe8473bae2b9dd73bbdef4bdef69fffffffffff"),
                (x"fffffffffffd084295c42108421084214a4210bfffffffffff"),
                (x"ffffffffffa10a5a50a408421084847508421094ffffffffff"),
                (x"fffffffdce2148ea50a4294a5294842d0a42048effffffffff"),
                (x"fffffffdce2148ea50a4294a5294842d0a42048effffffffff"),
                (x"fffffffc00710b4000a421084210842d1c4210b4a53fffffff"),
                (x"fffffffc004b1c0a508108421084212500421424003fffffff"),
                (x"ffffffffff03000738810842120421215c42058c003fffffff"),
                (x"fffffffffffffff73884f7bde2048473ba00312c003fffffff"),
                (x"fffffffffffffff73884f7bde2048473ba00312c003fffffff"),
                (x"fffffffffffffff003de6318c077bdef41ff8000ffffffffff"),
                (x"fffffffffffffffffc1d18c7d0018c603fffffffffffffffff"),
                (x"ffffffffffffffffffecefbcc0018c603fffffffffffffffff"),
                (x"fffffffffffffffffd8cb5acc0000007ffffffffffffffffff"),
                (x"fffffffffffffffffd8cb5acc0000007ffffffffffffffffff"),
                (x"fffffffffffffffffc0c6318c07fffffffffffffffffffffff"),

                -- 2_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffdce739d5ad6b5739dffffffffffffffff"),
                (x"fffffffffffffee73aa845ef7ba2b5aa2ae73bffffffffffff"),
                (x"fffffffffffffee73aa845ef7ba2b5aa2ae73bffffffffffff"),
                (x"ffffffffffffdd542117bdef7bdef7ba10845ebfffffffffff"),
                (x"fffffffffffbaa8ad508456b5ad508bdd15aa2eeffffffffff"),
                (x"ffffffffff7551542115aa108ba2b5aa2e8456f5ffffffffff"),
                (x"ffffffffff7551542115aa108ba2b5aa2e8456f5ffffffffff"),
                (x"ffffffffff756a8422a842117455294bab5ad5d573bfffffff"),
                (x"fffffffdcead508ad508aa108aa6f7bdd2e7393573bfffffff"),
                (x"fffffffdceaa11542115adee8adef7bdef7bdd3573bfffffff"),
                (x"ffffffbab5aa2b5422ae45ef54def7bdef7bdd2effffffffff"),
                (x"ffffffbab5455c8ad5ce45ef5bdef7bdef7bdd9dffffffffff"),
                (x"ffffffbab5455c8ad5ce45ef5bdef7bdef7bdd9dffffffffff"),
                (x"fffffed6b5455c8ad5ce42115ba58c632f7bdc1fffffffffff"),
                (x"fffffed5ceabab5739ceaa115ba4a5002f7bdc1fffffffffff"),
                (x"fffffed5ceabaaeef5d7aa10eba484002f7bdc1fffffffffff"),
                (x"fffffff5ce73abdef7a97210ebdc8439ef7bdc1fffffffffff"),
                (x"fffffff5ce73abdef7a97210ebdc8439ef7bdc1fffffffffff"),
                (x"fffffff5ceebabd73bb4756aebdc8491ef7bdc1fffffffffff"),
                (x"ffffffffbda75dd73bbd739c9bdef7bdef7bdc1fffffffffff"),
                (x"fffffffffffd3bd73bbda39c9bdef7bdef7ba41fffffffffff"),
                (x"ffffffffffffff4ef694a528c4def7bdee9483ffffffffffff"),
                (x"ffffffffffffff4ef694a528c4def7bdee9483ffffffffffff"),
                (x"fffffffffffffffffe94294b46318c6300007fffffffffffff"),
                (x"fffffffffffffffffe8520424210842fa9ffffffffffffffff"),
                (x"fffffffffffffffa50a520421290210fa9ffffffffffffffff"),
                (x"fffffffffffffffa50a521081214a52fbd4a7fffffffffffff"),
                (x"fffffffffffffffa50a521081214a52fbd4a7fffffffffffff"),
                (x"fffffffffffffffa50ae290852148427bd4a7fffffffffffff"),
                (x"ffffffffffffff4294b420421214840fbd4a7fffffffffffff"),
                (x"fffffffffffffee294b4a10810b8840fbd4a7fffffffffffff"),
                (x"ffffffffffffffd7389420421a50210fbd4a7fffffffffffff"),
                (x"ffffffffffffffd7389420421a50210fbd4a7fffffffffffff"),
                (x"ffffffffffffffdef7a475289bd0840f7bffffffffffffffff"),
                (x"fffffffffffffe0ef58ceb9ce213bdef7bffffffffffffffff"),
                (x"fffffffffffffe0633bde80000018c633fffffffffffffffff"),
                (x"fffffffffffffe06318c6001ff80006319ffffffffffffffff"),
                (x"fffffffffffffe06318c6001ff80006319ffffffffffffffff"),
                (x"fffffffffffffff0018cb3180fffffffffffffffffffffffff"),

                -- 2_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5ad5ce77fffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5ad5ce77fffffffffffff"),
                (x"ffffffffffffdd5ad6a8bdef5aa2f7ba115ab9dfffffffffff"),
                (x"fffffffffffbaa8bdef74211745ef7bdee8422aeffffffffff"),
                (x"fffffffffffd50842108bdee845ef7456a842115ffffffffff"),
                (x"fffffffffffd50842108bdee845ef7456a842115ffffffffff"),
                (x"ffffffffff756a8bdef742117422b5aa2f7ba11573bfffffff"),
                (x"ffffffffff756b5ad6a8bb9d545508bdd08456b573bfffffff"),
                (x"ffffffffbdad508ad5c9ba52eab929ba5d5aa2b5ad5dffffff"),
                (x"ffffffffbdaa11773937bdef7bdef7bdd2e7210ead5dffffff"),
                (x"fffffffdce456f573af7bdef7bdef7bdeee7550ead6aefffff"),
                (x"fffffffdce456f573af7bdef7bdef7bdeee7550ead6aefffff"),
                (x"fffffffdce43af573af7bdef7bdef7bdeee756ee73aaefffff"),
                (x"fffffff5ceaf50e4a58c65ef7bdef7631894bafd73aaeeffff"),
                (x"fffffff6b57250ebdca005ef7bdef7000b7bb909739d5effff"),
                (x"fffffff6b575eaebdc8005ef7bdef700097bbab773bb5effff"),
                (x"fffffff6b575eaebdc8005ef7bdef700097bbab773bb5effff"),
                (x"fffffff5ce702bdbdc873def7bdef739c97bf6a0ef40eeffff"),
                (x"ffffffffbd701c0bdc923def7bdef73c897b81c0ef41d07fff"),
                (x"ffffffffbde83a04a6f7bdef7bdef7bdee9483a0003e0fffff"),
                (x"ffffffffff0000063137bdef7bdef7bdd2c60000ffffffffff"),
                (x"ffffffffff0000063137bdef7bdef7bdd2c60000ffffffffff"),
                (x"ffffffffffffe850000c4a537bdd294b0052969fffffffffff"),
                (x"fffffffffffd0a5295c46318c6318c614842129fffffffffff"),
                (x"ffffffffff750a5294242109ef7884211c1090b4ffffffffff"),
                (x"fffffffe942908e000a10843ef78210b8a108494ffffffffff"),
                (x"fffffffe942908e000a10843ef78210b8a108494ffffffffff"),
                (x"fffffffdce214a5000a40843ef7821090a420424a53fffffff"),
                (x"fffffffe94611c0084052109ef78842140421024a53fffffff"),
                (x"fffffffc004b01f000a40909ef7884090042108e003fffffff"),
                (x"ffffffffff003ff000810909ef788421004239c5003fffffff"),
                (x"ffffffffff003ff000810909ef788421004239c5003fffffff"),
                (x"fffffffffffffff001c42109def7bd23800026e0ffffffffff"),
                (x"fffffffffffffffffc0eafbdeef7bdef7fff801fffffffffff"),
                (x"ffffffffffffffffffe0e8c7ee818c67ffffffffffffffffff"),
                (x"ffffffffffffffffffe067bdd6000007ffffffffffffffffff"),
                (x"ffffffffffffffffffe067bdd6000007ffffffffffffffffff"),
                (x"ffffffffffffffffffe065ad6603ffffffffffffffffffffff"),

                -- 2_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff739cead6b5ab9ce73bfffffffffffffffff"),
                (x"ffffffffffffdcead515aa117bdd08455ce77fffffffffffff"),
                (x"ffffffffffffdcead515aa117bdd08455ce77fffffffffffff"),
                (x"fffffffffffd6e842117bdef7bdef7ba115abbffffffffffff"),
                (x"ffffffffff75d15422f7456b5ad508422a8455dfffffffffff"),
                (x"ffffffffffadea8bdd15aa117422b5aa115aa2aeffffffffff"),
                (x"ffffffffffadea8bdd15aa117422b5aa115aa2aeffffffffff"),
                (x"fffffffdceabab5ad5c94d6a8ba10845508456aeffffffffff"),
                (x"fffffffdceaa5ce4a6f7ba535422b5422a8422b573bfffffff"),
                (x"fffffffdceaa6f7bdef7bdef545eb5aa115aa11573bfffffff"),
                (x"ffffffffff726f7bdef7bdee9add0875515ad515ad5dffffff"),
                (x"ffffffffffeb2f7bdef7bdef7add0873aa843aa8ad5dffffff"),
                (x"ffffffffffeb2f7bdef7bdef7add0873aa843aa8ad5dffffff"),
                (x"fffffffffff82f7bdd8c62537aa10873aa843aa8ad6bdfffff"),
                (x"fffffffffff82f7bdc002a537aa2b5739d5ad5d573abdfffff"),
                (x"fffffffffff82f7bdc0022537722b5bbbae755d573abdfffff"),
                (x"fffffffffff82f7bdce725ef7721ce4f7bded5ce73bbffffff"),
                (x"fffffffffff82f7bdce725ef7721ce4f7bded5ce73bbffffff"),
                (x"fffffffffff82f7bdcf225ef7755cea75dded5dd73bbffffff"),
                (x"fffffffffff82f7bdef7bdef74b9ceef5ddebbb4ef7fffffff"),
                (x"fffffffffff8137bdef7bdef74ba94ef5ddef69fffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a53b4a7fffffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a53b4a7fffffffffffff"),
                (x"fffffffffffffe00018c6318ca14a5a53fffffffffffffffff"),
                (x"fffffffffffffffa53c521084204842d3fffffffffffffffff"),
                (x"fffffffffffffffa53c109085084842969ffffffffffffffff"),
                (x"ffffffffffffff4f7bc5294a4090842969ffffffffffffffff"),
                (x"ffffffffffffff4f7bc5294a4090842969ffffffffffffffff"),
                (x"ffffffffffffff4f7bc4214a4290a57169ffffffffffffffff"),
                (x"ffffffffffffff4f7bc1214a408484a14b4a7fffffffffffff"),
                (x"ffffffffffffff4f7bc1239c109294a14ae77fffffffffffff"),
                (x"ffffffffffffff4f7bc10d29408484a11ddeffffffffffffff"),
                (x"ffffffffffffff4f7bc10d29408484a11ddeffffffffffffff"),
                (x"fffffffffffffffef7a1252974d1ce277bdeffffffffffffff"),
                (x"fffffffffffffffef7bded6b573bbd633a007fffffffffffff"),
                (x"fffffffffffffffffd8c60000003bdef58007fffffffffffff"),
                (x"fffffffffffffff6318c0001ff818c6318007fffffffffffff"),
                (x"fffffffffffffff6318c0001ff818c6318007fffffffffffff"),
                (x"fffffffffffffffffffffffff032d66301ffffffffffffffff"),

                -- 2_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce73bfffffffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5756ae77fffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5756ae77fffffffffffff"),
                (x"ffffffffffffdd5ad517ad6a8aa2b5aa115ad5dfffffffffff"),
                (x"fffffffffffbaa8422a8bd6b7422b5422b5aa2aeffffffffff"),
                (x"fffffffffffd51742115ba117455084550842115ffffffffff"),
                (x"fffffffffffd51742115ba117455084550842115ffffffffff"),
                (x"ffffffffff722f742108421084550842108422f573bfffffff"),
                (x"ffffffffff75ef7bdd084211742108ba10845d1573bfffffff"),
                (x"ffffffffbdadee8422f7ba117ba2f7bdef7ba2b5ad7bffffff"),
                (x"ffffffffbd45d0842108bdef7bdef7bdd0842115ad7bffffff"),
                (x"fffffff5ce42108421084211742108ba10842115ad7bffffff"),
                (x"fffffff5ce42108421084211742108ba10842115ad7bffffff"),
                (x"fffffff6b5455084210842108421084550842115ad5dffffff"),
                (x"fffffeb9084550842108421084210845508422a8ad5ddfffff"),
                (x"fffff75508aa115422a8421084210845508422a8ad5ddfffff"),
                (x"fffff75508722a8422a84210842108ad515aa1c8739ddfffff"),
                (x"fffff75508722a8422a84210842108ad515aa1c8739ddfffff"),
                (x"fffffeb908756a8421c8aa1154210875515ad5d5739ddfffff"),
                (x"fffffff6b5ed5c8ad7a8aa10e422b575515abab573bbffffff"),
                (x"fffffffc00ef5c873bb57210e422b573ab5abaae73bbffffff"),
                (x"fffffffffffffbd297aeed6bdad5ceebaae775ceef7fffffff"),
                (x"fffffffffffffbd297aeed6bdad5ceebaae775ceef7fffffff"),
                (x"ffffffffffffe85210bdef7a5777bd2f5dde93bdffffffffff"),
                (x"ffffffffffffca4210a52108421084211c529094ffffffffff"),
                (x"fffffffffffd08421094710810842109094a14a4a53fffffff"),
                (x"fffffffffffb881210b429085294a5290b4a3885211dffffff"),
                (x"fffffffffffb881210b429085294a5290b4a3885211dffffff"),
                (x"ffffffffffa50a4211d42908421084210a0050a47381ffffff"),
                (x"ffffffffff0102521014210810842109094a01ccf781ffffff"),
                (x"ffffffffff03181211c520421084210848e7000c003fffffff"),
                (x"ffffffffff0312c003ae7108127bdef108e77fffffffffffff"),
                (x"ffffffffff0312c003ae7108127bdef108e77fffffffffffff"),
                (x"fffffffffff8000ffc1def7bd0318c67bc007fffffffffffff"),
                (x"ffffffffffffffffffe063180074631f41ffffffffffffffff"),
                (x"ffffffffffffffffffe063180033deeb3fffffffffffffffff"),
                (x"ffffffffffffffffffff00000032d6b319ffffffffffffffff"),
                (x"ffffffffffffffffffff00000032d6b319ffffffffffffffff"),
                (x"fffffffffffffffffffffffff0318c6301ffffffffffffffff"),

                -- 2_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffdce739d5ad6b5739dffffffffffffffff"),
                (x"fffffffffffffee73aa845ef7ba2b5aa2ae73bffffffffffff"),
                (x"fffffffffffffee73aa845ef7ba2b5aa2ae73bffffffffffff"),
                (x"ffffffffffffdd542117bdef7bdef7ba10845ebfffffffffff"),
                (x"fffffffffffbaa8ad508456b5ad508bdd15aa2eeffffffffff"),
                (x"ffffffffff7551542115aa108ba2b5aa2e8456f5ffffffffff"),
                (x"ffffffffff7551542115aa108ba2b5aa2e8456f5ffffffffff"),
                (x"ffffffffff756a8422a842117455294bab5ad5d573bfffffff"),
                (x"ffffffffff756a842108aa108aa6f7bdd2e7393573bfffffff"),
                (x"fffffffdcead6a8ad508adee8adef7bdef7bdd3573bfffffff"),
                (x"fffffffdcead508ad51545ef54def7bdef7bdd2effffffffff"),
                (x"fffffffdceab908ad51545ef5bdef7bdef7bdd9dffffffffff"),
                (x"fffffffdceab908ad51545ef5bdef7bdef7bdd9dffffffffff"),
                (x"fffffffdceab9157390e42115ba58c632f7bdc1fffffffffff"),
                (x"ffffffffbdab91573aaeaa115ba4a5002f7bdc1fffffffffff"),
                (x"ffffffffbdab915739d7aa10eba484002f7bdc1fffffffffff"),
                (x"ffffffffbd776b5739c97210ebdc8439ef7bdc1fffffffffff"),
                (x"ffffffffbd776b5739c97210ebdc8439ef7bdc1fffffffffff"),
                (x"ffffffffbd776b5739d4756aebdc8491ef7bdc1fffffffffff"),
                (x"ffffffffffef5d5ef5dd739c9bdef7bdef7bdc1fffffffffff"),
                (x"fffffffffffd3aeef5dda39c9bdef7bdef7ba41fffffffffff"),
                (x"ffffffffffffff4ef694a528c4def7bdee9483ffffffffffff"),
                (x"ffffffffffffff4ef694a528c4def7bdee9483ffffffffffff"),
                (x"fffffffffffffffa50a5a39c56318c6300007fffffffffffff"),
                (x"ffffffffffffff4294812908525294a51c4253ffffffffffff"),
                (x"ffffffffffffff421081214a409484a78252d3ffffffffffff"),
                (x"fffffffffffffee29484214a4085cea7a852969fffffffffff"),
                (x"fffffffffffffee29484214a4085cea7a852969fffffffffff"),
                (x"ffffffffffffe852102ea1081091cea7a852ba9fffffffffff"),
                (x"ffffffffffffe8e294a50108421484a7bd4a149fffffffffff"),
                (x"ffffffffffffe942102e0108109421a7bd4a101fffffffffff"),
                (x"ffffffffffffc0c6318071084084a5efbd4a5c1fffffffffff"),
                (x"ffffffffffffc0c6318071084084a5efbd4a5c1fffffffffff"),
                (x"fffffffffffffe04a6e0ed6b5efbdef7400003ffffffffffff"),
                (x"fffffffffffffe00001def7bdef7bdef41ffffffffffffffff"),
                (x"fffffffffffffe06318000000ef863603fffffffffffffffff"),
                (x"fffffffffffffe06318c07fe0677de6301ffffffffffffffff"),
                (x"fffffffffffffe06318c07fe0677de6301ffffffffffffffff"),
                (x"fffffffffffffffffffffffff032d6b301ffffffffffffffff"),

                -- 2_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffee739ce739ce77ffffffffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5ad5ce77fffffffffffff"),
                (x"fffffffffffffffad6b5ad6b5756b5ad5ce77fffffffffffff"),
                (x"ffffffffffffdd5ad6a8bdef5aa2f7ba115ab9dfffffffffff"),
                (x"fffffffffffbaa8bdef74211745ef7bdee8422aeffffffffff"),
                (x"fffffffffffd50842108bdee845ef7456a842115ffffffffff"),
                (x"fffffffffffd50842108bdee845ef7456a842115ffffffffff"),
                (x"ffffffffff756a8bdef742117422b5aa2f7ba11573bfffffff"),
                (x"ffffffffff756b5ad6a8bb9d545508bdd08456b573bfffffff"),
                (x"ffffffffbdad508ad5c9ba52eab929ba5d5aa2b573bbffffff"),
                (x"ffffffffbdaa11773937bdef7bdef7bdd2e72115ad7bffffff"),
                (x"ffffffbab5ab91573af7bdef7bdef7bdeee756f5ad5dffffff"),
                (x"ffffffbab5ab91573af7bdef7bdef7bdeee756f5ad5dffffff"),
                (x"ffffffbab573af573af7bdef7bdef7bdeee756eead5ddfffff"),
                (x"fffffebab5776ee4a58c65ef7bdef7631894b91dad5ddfffff"),
                (x"fffffed5ce7250ebdca005ef7bdef7000b7bb909739ddfffff"),
                (x"fffffed7bd75eaebdc8005ef7bdef700097bbab7ef5ddfffff"),
                (x"fffffed7bd75eaebdc8005ef7bdef700097bbab7ef5ddfffff"),
                (x"fffffebbbde82bdbdc873def7bdef739c97bf6a073bbffffff"),
                (x"fffff07400e81c0bdc923def7bdef73c897b81c073bbffffff"),
                (x"ffffff83ffe83a04a6f7bdef7bdef7bdee9483a0ef7fffffff"),
                (x"ffffffffff07c0063137bdef7bdef7bdd2c60000ffffffffff"),
                (x"ffffffffff07c0063137bdef7bdef7bdd2c60000ffffffffff"),
                (x"ffffffffffffe852940c4a537bdd294b0000169fffffffffff"),
                (x"ffffffffffffe84210856318c6318c611c5294b4ffffffffff"),
                (x"fffffffffffd0a4085c12109ef788421025294b473bfffffff"),
                (x"fffffffffffd081084ae0843ef7821084a0038842969ffffff"),
                (x"fffffffffffd081084ae0843ef7821084a0038842969ffffff"),
                (x"ffffffffffa1021210a40843ef7821090a0014a5211dffffff"),
                (x"ffffffffffa1024210052109ef788421401081c46329ffffff"),
                (x"ffffffffff03884210040909ef7884090a007c0c4a41ffffff"),
                (x"ffffffffff015ce210042109ef78840848007fe0003fffffff"),
                (x"ffffffffff015ce210042109ef78840848007fe0003fffffff"),
                (x"fffffffffff82e90000e277bdef484211c007fffffffffffff"),
                (x"ffffffffffffc00ffffdef7bdf7bdeab81ffffffffffffffff"),
                (x"ffffffffffffffffffff63180ef863e83fffffffffffffffff"),
                (x"ffffffffffffffffffff00000677de603fffffffffffffffff"),
                (x"ffffffffffffffffffff00000677de603fffffffffffffffff"),
                (x"fffffffffffffffffffffffe065ad6603fffffffffffffffff"),

                -- 2_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff739cead6b5ab9ce73bfffffffffffffffff"),
                (x"ffffffffffffdcead515aa117bdd08455ce77fffffffffffff"),
                (x"ffffffffffffdcead515aa117bdd08455ce77fffffffffffff"),
                (x"fffffffffffd6e842117bdef7bdef7ba115abbffffffffffff"),
                (x"ffffffffff75d15422f7456b5ad508422a8455dfffffffffff"),
                (x"ffffffffffadea8bdd15aa117422b5aa115aa2aeffffffffff"),
                (x"ffffffffffadea8bdd15aa117422b5aa115aa2aeffffffffff"),
                (x"fffffffdceabab5ad5c94d6a8ba10845508456aeffffffffff"),
                (x"fffffffdceaa5ce4a6f7ba535422b542108456aeffffffffff"),
                (x"fffffffdceaa6f7bdef7bdef545eb5422a8456b573bfffffff"),
                (x"ffffffffff726f7bdef7bdee9add08aa2a8422b573bfffffff"),
                (x"ffffffffffeb2f7bdef7bdef7add08aa2a8421d573bfffffff"),
                (x"ffffffffffeb2f7bdef7bdef7add08aa2a8421d573bfffffff"),
                (x"fffffffffff82f7bdd8c62537aa108721d5aa1d573bfffffff"),
                (x"fffffffffff82f7bdc002a537aa2b5755d5aa1d5ef7fffffff"),
                (x"fffffffffff82f7bdc0022537722b5bb9d5aa1d5ef7fffffff"),
                (x"fffffffffff82f7bdce725ef7721ce4b9d5ad7aeef7fffffff"),
                (x"fffffffffff82f7bdce725ef7721ce4b9d5ad7aeef7fffffff"),
                (x"fffffffffff82f7bdcf225ef7755cea39d5ad7aeef7fffffff"),
                (x"fffffffffff82f7bdef7bdef74b9ceebbb5abbbdffffffffff"),
                (x"fffffffffff8137bdef7bdef74ba94ebbae7769fffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a53b4a7fffffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a53b4a7fffffffffffff"),
                (x"fffffffffffffe00018c6318c2ba942969ffffffffffffffff"),
                (x"ffffffffffffe8473a94a5284290a5090b4a7fffffffffffff"),
                (x"ffffffffffffe85087d4214a12148409094a7fffffffffffff"),
                (x"fffffffffffd0a5a53d47042121484210ae77fffffffffffff"),
                (x"fffffffffffd0a5a53d47042121484210ae77fffffffffffff"),
                (x"fffffffffffd1c5a53d47108109294704852d3ffffffffffff"),
                (x"fffffffffff90b4f7bd4214a421000294ae753ffffffffffff"),
                (x"fffffffffff8094f7bd4094a10900070494a53ffffffffffff"),
                (x"fffffffffff82f4f7bdd28421211ce0318c603ffffffffffff"),
                (x"fffffffffff82f4f7bdd28421211ce0318c603ffffffffffff"),
                (x"ffffffffffffc00003bef7bdd213bd05d2007fffffffffffff"),
                (x"fffffffffffffff003bdef7bdef7bde800007fffffffffffff"),
                (x"fffffffffffffffffc0c1fbdd000000318007fffffffffffff"),
                (x"fffffffffffffff0018cf77ac07c006318007fffffffffffff"),
                (x"fffffffffffffff0018cf77ac07c006318007fffffffffffff"),
                (x"fffffffffffffff00196b3180fffffffffffffffffffffffff"),

                -- 3_character_0_0
                (x"fffffffffffffffffffef7bdef7bdef7bfffffffffffffffff"),
                (x"ffffffffffffffff7bc739ce739ce739fdef7fffffffffffff"),
                (x"ffffffffffffffe39ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffffe39ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffe8718c6318c6318c6318ce739e9fffffffffff"),
                (x"fffffffffffd3c318c6318c6318c6318c6739fd4ffffffffff"),
                (x"fffffffffffd0e318c6318c6318c6318c6739cf4ffffffffff"),
                (x"fffffffffffd0e318c6318c6318c6318c6739cf4ffffffffff"),
                (x"ffffffffffa786318ce318c6318c6318ce739cfea53fffffff"),
                (x"ffffffffffa1c6318ce718c6318c6319ce739cfea53fffffff"),
                (x"ffffffffffa0ce318ce739ce739ce739ce739cfea53fffffff"),
                (x"ffffffffffa0fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa1fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa1fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa7bc718c7e39ce739ce73f8e739fdea53fffffff"),
                (x"ffffffffffa7bde39c7e39ce739ce7f78e73fbdea53fffffff"),
                (x"fffffffffffd3de39ce7f1ce739ce7f1ce73fbd4a53fffffff"),
                (x"fffffffffffd3def78e7f7bc739fdef1cfef7bd4ffffffffff"),
                (x"fffffffffffd3def78e7f7bc739fdef1cfef7bd4ffffffffff"),
                (x"ffffffffffffe9ef7bc73d29ef7a9439fdef7a9fffffffffff"),
                (x"ffffffffffffff4f7bdef5294a7a94f7bdef53ffffffffffff"),
                (x"ffffffffffffe87a529e3fbc719fde3fa94a1e9fffffffffff"),
                (x"fffffffffffd0e3f7a9df77b4a52940529ef0cf4ffffffffff"),
                (x"fffffffffffd0e3f7a9df77b4a52940529ef0cf4ffffffffff"),
                (x"ffffffffffa7867f7a9df7bdef7bdef77bef1c7ea53fffffff"),
                (x"fffffffe94a78fef7a9df7bdef7bdef7a9ef78fea529ffffff"),
                (x"fffffffe94f5294f7a94efbd4f53def769ef5294f7a9ffffff"),
                (x"ffffffffbda7bd400294a529def694a5280053dea53bffffff"),
                (x"ffffffffbda7bd400294a529def694a5280053dea53bffffff"),
                (x"fffffffe94ed00000294ef7bdef7bded28000014ef69ffffff"),
                (x"fffffffe94a52940029e38c67f1c633fa8005294a529ffffff"),
                (x"ffffffffffa528000294f1cfea78e7f528000294a53fffffff"),
                (x"fffffffffffffffa53c7a528000294a1fd4a7fffffffffffff"),
                (x"fffffffffffffffa53c7a528000294a1fd4a7fffffffffffff"),
                (x"fffffffffffffffa529e19cfea78e71fa94a7fffffffffffff"),
                (x"fffffffffffffff00294a529405294a528007fffffffffffff"),
                (x"fffffffffffffffffc1ef529405294f781ffffffffffffffff"),
                (x"fffffffffffffffffc14f5280f8294f501ffffffffffffffff"),
                (x"fffffffffffffffffc14f5280f8294f501ffffffffffffffff"),
                (x"fffffffffffffffffc1e3fbc0f83de3f81ffffffffffffffff"),

                -- 3_character_0_1
                (x"fffffffffffffffffe94a5294f7bdef7bfffffffffffffffff"),
                (x"ffffffffffffff4a53de38c6318c6339fdef7fffffffffffff"),
                (x"ffffffffffffe9e39ce739ce738c6318c673fbffffffffffff"),
                (x"ffffffffffffe9e39ce739ce738c6318c673fbffffffffffff"),
                (x"fffffffffffd3c739ce739ce318c631f9e31bfdfffffffffff"),
                (x"fffffffffffd0e739ce718c6318c63f0c65295ffffffffffff"),
                (x"ffffffffffa78e7f78e319cfef1fde1bfc31d0b4ffffffffff"),
                (x"ffffffffffa78e7f78e319cfef1fde1bfc31d0b4ffffffffff"),
                (x"ffffffffffa78fef78e7f7bc7f78637f803180b4ffffffffff"),
                (x"fffffffe94f7bde39cfef529418fdef500f78074ffffffffff"),
                (x"fffffffe94f7bde39fd4a3de37fbdef500f781f4ffffffffff"),
                (x"fffffffe94f7bdef780f7fbdef7bdef7a9ef51e0ffffffffff"),
                (x"fffffffe94f7bdea501ef7bdef5000003def781fffffffffff"),
                (x"fffffffe94f7bdea501ef7bdef5000003def781fffffffffff"),
                (x"ffffffffffa7bdef7814f7bdea0339000000001fffffffffff"),
                (x"ffffffffffa7bd4f7bd405294a0339ce4e739c1fffffffffff"),
                (x"fffffffffffd3d4f7a9405294783399cce739c1fffffffffff"),
                (x"fffffffffffd294a529405294f3fde9d0652947fffffffffff"),
                (x"fffffffffffd294a529405294f3fde9d0652947fffffffffff"),
                (x"fffffffffffffd4a529405294f79efa0def780b4ffffffffff"),
                (x"ffffffffffffff4a529405294f7bdea3c0f78074ffffffffff"),
                (x"fffffffffffffffffe94a0014a7bdea3e8f7801fffffffffff"),
                (x"fffffffffffffffffc14a528000294a5280003ffffffffffff"),
                (x"fffffffffffffffffc14a528000294a5280003ffffffffffff"),
                (x"fffffffffffffff003c7a529da5294a501ffffffffffffffff"),
                (x"fffffffffffffffa5063f529df77de3fa9ffffffffffffffff"),
                (x"fffffffffffffe0f78fe38c67a50e739fdffffffffffffffff"),
                (x"fffffffffffffe0f7a871f7b400294f7a9ffffffffffffffff"),
                (x"fffffffffffffe0f7a871f7b400294f7a9ffffffffffffffff"),
                (x"fffffffffffffe0a5287ed29e1f800a501ffffffffffffffff"),
                (x"fffffffffffffff0029eed2873f800ed01ffffffffffffffff"),
                (x"fffffffffffffff00014a529ef500019e9ffffffffffffffff"),
                (x"fffffffffffffff00280a5294003de3d29ffffffffffffffff"),
                (x"fffffffffffffff00280a5294003de3d29ffffffffffffffff"),
                (x"fffffffffffffffffc1400000a5294f53fffffffffffffffff"),
                (x"ffffffffffffffffffe0a7bc719fdea7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0a7bdef529407ffffffffffffffffff"),
                (x"ffffffffffffffffffffa5294a5000ffffffffffffffffffff"),
                (x"ffffffffffffffffffffa5294a5000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bde3f800ffffffffffffffffffff"),

                -- 3_character_0_2
                (x"fffffffffffffffffffff7bdea5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffdef1ce739ce7f7a94a7fffffffffffff"),
                (x"ffffffffffffff4f78e718c6318c6318cfef53ffffffffffff"),
                (x"ffffffffffffff4f78e718c6318c6318cfef53ffffffffffff"),
                (x"ffffffffffffe9e39c6318c6318c6318c673fa9fffffffffff"),
                (x"fffffffffffd3c718c6339cfef78e739c6319fd4ffffffffff"),
                (x"fffffffffffd0e339ce7f3de5295eff7bc739fd4ffffffffff"),
                (x"fffffffffffd0e339ce7f3de5295eff7bc739fd4ffffffffff"),
                (x"ffffffffffa786739cef294a3a78a51bfdef7bdea53fffffff"),
                (x"ffffffffffa787e39de57d28307a9478dfef7a9ea53fffffff"),
                (x"ffffffffffa1fc77bcaf18003078007f86f7fa9ea53fffffff"),
                (x"ffffffffffa1e9e295e318003a78007fbc31fa94a53fffffff"),
                (x"ffffffffffa01efa53cf1d283a7a947fbd4a3de0a53fffffff"),
                (x"ffffffffffa01efa53cf1d283a7a947fbd4a3de0a53fffffff"),
                (x"ffffffffffa03de0001e78c637f9eff780007bc0a53fffffff"),
                (x"ffffffffffa529e0032005294a52940032007a94a53fffffff"),
                (x"ffffffffffa501400339c9ce739ce7ce72005014a53fffffff"),
                (x"fffffffffff8014a53339fbd4a53de9cf34a5000ffffffffff"),
                (x"fffffffffff8014a53339fbd4a53de9cf34a5000ffffffffff"),
                (x"ffffffffffffc1ea5333f14a529463f4f34a781fffffffffff"),
                (x"ffffffffffffc14f787428c63079ef1d1fef501fffffffffff"),
                (x"fffffffffffd3d4f79f47800307800f51fef53d4ffffffffff"),
                (x"fffffffe94a7867a53d47d28307a94f53d4a1c7ea529ffffff"),
                (x"fffffffe94a7867a53d47d28307a94f53d4a1c7ea529ffffff"),
                (x"ffffffd0e719cfea5294a3deff7bdea5294a78e718cf4fffff"),
                (x"fffffa1fdea5294a529df5294a5294f7694a5294a53c7a7fff"),
                (x"fffffa1e94ef694a53dd39ce739ce73f7d4a529def687a7fff"),
                (x"fffff053bda529400294f7bdef7bdef528005294a53b407fff"),
                (x"fffff053bda529400294f7bdef7bdef528005294a53b407fff"),
                (x"ffffff8294a0cf400294a5294a5294a5280050e3a5280fffff"),
                (x"fffffffc00f1cf400294a77bdef7bda5280050e7f7800fffff"),
                (x"fffffffc00a7bc000294f1ce318ce7f5280003dea501ffffff"),
                (x"ffffffffff0001f00014a7bc739fdea500007c00003fffffff"),
                (x"ffffffffff0001f00014a7bc739fdea500007c00003fffffff"),
                (x"fffffffffffffffa53c7a529405294a1fd4a7fffffffffffff"),
                (x"fffffffffffffff0029e19cf4050e71fa8007fffffffffffff"),
                (x"fffffffffffffff00294a528000294a528007fffffffffffff"),
                (x"fffffffffffffffffc1e1fbc0f83de1f81ffffffffffffffff"),
                (x"fffffffffffffffffc1e1fbc0f83de1f81ffffffffffffffff"),
                (x"fffffffffffffffffc14a5280f8294a501ffffffffffffffff"),

                -- 3_character_0_3
                (x"ffffffffffffffffffdef7bdea5294a53fffffffffffffffff"),
                (x"ffffffffffffffef78e718c6318ce7f7a94a7fffffffffffff"),
                (x"fffffffffffffc718c6318c6739ce739cfef53ffffffffffff"),
                (x"fffffffffffffc718c6318c6739ce739cfef53ffffffffffff"),
                (x"ffffffffffff9e37bfc318c6319ce739ce73fa9fffffffffff"),
                (x"fffffffffffbca518c7e18c6318c6339ce739e9fffffffffff"),
                (x"ffffffffffa1683f79e3f1cfef1c6319fc739fd4ffffffffff"),
                (x"ffffffffffa1683f79e3f1cfef1c6319fc739fd4ffffffffff"),
                (x"ffffffffffa1403003cf1fbde3fbde39fdef1fd4ffffffffff"),
                (x"ffffffffffa0c0f0029ef0c63a53def1cfef7bdea53fffffff"),
                (x"ffffffffffa3c0f0029ef7bcf1be94a78fef7bdea53fffffff"),
                (x"ffffffffff03e9ea53def7bdef79ef783def7bdea53fffffff"),
                (x"fffffffffff83def78000529ef7bdef029ef7bdea53fffffff"),
                (x"fffffffffff83def78000529ef7bdef029ef7bdea53fffffff"),
                (x"fffffffffff800000000c8014f7bdea03def7bd4ffffffffff"),
                (x"fffffffffff80e739f39c8014a5000a7bd4a7bd4ffffffffff"),
                (x"fffffffffff80e739e73c800fa5000a53d4a7a9fffffffffff"),
                (x"fffffffffff8ca518e93f3dfea5000a5294a529fffffffffff"),
                (x"fffffffffff8ca518e93f3dfea5000a5294a529fffffffffff"),
                (x"ffffffffffa140f7bc747fbdea5000a5294a7bffffffffffff"),
                (x"ffffffffffa0c0f001f4f7bdea5000a529ffffffffffffffff"),
                (x"fffffffffff800fa51f4f7bd4a0294a53fffffffffffffffff"),
                (x"ffffffffffffc00a5294a000005294a03fffffffffffffffff"),
                (x"ffffffffffffc00a5294a000005294a03fffffffffffffffff"),
                (x"fffffffffffffff00294a5294ed2943f81ffffffffffffffff"),
                (x"fffffffffffffffa53c7f77beed3de18e9ffffffffffffffff"),
                (x"ffffffffffffffff78e73d29438ce7f1fc007fffffffffffff"),
                (x"fffffffffffffffa53dea0000a74633d3c007fffffffffffff"),
                (x"fffffffffffffffa53dea0000a74633d3c007fffffffffffff"),
                (x"fffffffffffffff0029407bc3f53bd3d28007fffffffffffff"),
                (x"fffffffffffffff0029d07bc73d3bdf501ffffffffffffffff"),
                (x"fffffffffffffffa50e30529ef5294a001ffffffffffffffff"),
                (x"fffffffffffffffa5287f0000a52940501ffffffffffffffff"),
                (x"fffffffffffffffa5287f0000a52940501ffffffffffffffff"),
                (x"fffffffffffffffffe9ea529400000a03fffffffffffffffff"),
                (x"fffffffffffffffffff4f1ce33fa9407ffffffffffffffffff"),
                (x"ffffffffffffffffffe0a529ef7a9407ffffffffffffffffff"),
                (x"ffffffffffffffffffff05294a5294ffffffffffffffffffff"),
                (x"ffffffffffffffffffff05294a5294ffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc7f7800ffffffffffffffffffff"),

                -- 3_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffef7bdef7bdef7bfffffffffffffffff"),
                (x"ffffffffffffffff7bc739ce739ce739fdef7fffffffffffff"),
                (x"ffffffffffffffff7bc739ce739ce739fdef7fffffffffffff"),
                (x"ffffffffffffffe39ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffe8718c6318c6318c6318ce739e9fffffffffff"),
                (x"fffffffffffd3c318c6318c6318c6318c6739fd4ffffffffff"),
                (x"fffffffffffd3c318c6318c6318c6318c6739fd4ffffffffff"),
                (x"fffffffffffd0e318c6318c6318c6318c6739cf4ffffffffff"),
                (x"ffffffffffa786318ce318c6318c6318ce739cfea53fffffff"),
                (x"ffffffffffa1c6318ce718c6318c6319ce739cfea53fffffff"),
                (x"ffffffffffa0ce318ce739ce739ce739ce739cfea53fffffff"),
                (x"ffffffffffa0fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa0fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa1fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa7bc718c7e39ce739ce73f8e739fdea53fffffff"),
                (x"ffffffffffa7bde39c7e39ce739ce7f78e73fbdea53fffffff"),
                (x"fffffffffffd3de39ce7f1ce739ce7f1ce73fbd4a53fffffff"),
                (x"fffffffffffd3de39ce7f1ce739ce7f1ce73fbd4a53fffffff"),
                (x"fffffffffffd3def78e7f7bc739fdef1cfef7bd4ffffffffff"),
                (x"ffffffffffffe9ef7bc73d29ef7a9439fdef7a9fffffffffff"),
                (x"ffffffffffffff4f7bdef5294a7a94f7bdef53ffffffffffff"),
                (x"ffffffffffffe9ea529df77b4a529405294a53ffffffffffff"),
                (x"ffffffffffffe9ea529df77b4a529405294a53ffffffffffff"),
                (x"fffffffffffd3c7f7a9df7bde1fbdef77bef7a9fffffffffff"),
                (x"ffffffffffa78fef7a9df7bdef7bdef7a9ef1e9fffffffffff"),
                (x"fffffffe94a53d4f7a94efbd4f7bdef769ef7a94ffffffffff"),
                (x"fffffffe94a7bd4f7a94a529def694a529ef5294a53fffffff"),
                (x"fffffffe94a7bd4f7a94a529def694a529ef5294a53fffffff"),
                (x"ffffffffffa5280003d4a5294a5294a03d4a53d4a53fffffff"),
                (x"ffffffffffa53b4a5294ef7bded294a03def7bb4003fffffff"),
                (x"fffffffffffd294003c719cfea78e7f529def694ffffffffff"),
                (x"ffffffffffffc000029ef5280053dea5014a5280ffffffffff"),
                (x"ffffffffffffc000029ef5280053dea5014a5280ffffffffff"),
                (x"fffffffffffffffffc1439cfe05294a5000003ffffffffffff"),
                (x"fffffffffffffffffc1ef5294f0294a03fffffffffffffffff"),
                (x"ffffffffffffffffffe0a1ce7f000007ffffffffffffffffff"),
                (x"ffffffffffffffffffff07bd4a03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bd4a03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff05294a03ffffffffffffffffffffff"),

                -- 3_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294f7bdef7bfffffffffffffffff"),
                (x"ffffffffffffff4a53de38c6318c6339fdef7fffffffffffff"),
                (x"ffffffffffffff4a53de38c6318c6339fdef7fffffffffffff"),
                (x"ffffffffffffe9e39ce739ce738c6318c673fbffffffffffff"),
                (x"fffffffffffd3c739ce739ce318c631f9e31bfdfffffffffff"),
                (x"fffffffffffd0e739ce718c6318c63f0c65295ffffffffffff"),
                (x"fffffffffffd0e739ce718c6318c63f0c65295ffffffffffff"),
                (x"ffffffffffa78e7f78e319cfef1fde1bfc31d0b4ffffffffff"),
                (x"ffffffffffa78fef78e7f7bc7f78637f803180b4ffffffffff"),
                (x"fffffffe94f7bde39cfef529418fdef500f78074ffffffffff"),
                (x"fffffffe94f7bde39fd4a3de37fbdef500f781f4ffffffffff"),
                (x"fffffffe94f7bdef780f7fbdef7bdef7a9ef51e0ffffffffff"),
                (x"fffffffe94f7bdef780f7fbdef7bdef7a9ef51e0ffffffffff"),
                (x"fffffffe94f7bdea501ef7bdef5000003def781fffffffffff"),
                (x"ffffffffffa7bdef7814f7bdea0339000000001fffffffffff"),
                (x"ffffffffffa7bd4f7bd405294a0339ce4e739c1fffffffffff"),
                (x"fffffffffffd3d4f7a9405294783399cce739c1fffffffffff"),
                (x"fffffffffffd3d4f7a9405294783399cce739c1fffffffffff"),
                (x"fffffffffffd294a529405294f3fde9d0652947fffffffffff"),
                (x"fffffffffffffd4a529405294f79efa0def780b4ffffffffff"),
                (x"fffffffffffffffa529405294f7bdea3c0f78074ffffffffff"),
                (x"fffffffffffffffffe94a0014a7bdea3e8f7801fffffffffff"),
                (x"fffffffffffffffffe94a0014a7bdea3e8f7801fffffffffff"),
                (x"fffffffffffffffffc14a77a000294a5280003ffffffffffff"),
                (x"fffffffffffffffffc1e3d29df5294a529ffffffffffffffff"),
                (x"fffffffffffffff003c31fbd4a77de3fa9ffffffffffffffff"),
                (x"fffffffffffffff003c7f5287a529439e9ffffffffffffffff"),
                (x"fffffffffffffff003c7f5287a529439e9ffffffffffffffff"),
                (x"fffffffffffffff0029ea1cfee9fdea7a9ffffffffffffffff"),
                (x"fffffffffffffe0a5014a7bd4e8c633fa9ffffffffffffffff"),
                (x"fffffffffffffe0f7a80a7bdda1c63f53fffffffffffffffff"),
                (x"ffffffffffffff4f7a9405294a0000053fffffffffffffffff"),
                (x"ffffffffffffff4f7a9405294a0000053fffffffffffffffff"),
                (x"fffffffffffffe0a53c7a000000294a53fffffffffffffffff"),
                (x"fffffffffffffe0a529e39cf4053de3fbfffffffffffffffff"),
                (x"fffffffffffffffa5294a5280a5294f53fffffffffffffffff"),
                (x"ffffffffffffffff7bd40001ffd3de3fa9ffffffffffffffff"),
                (x"ffffffffffffffff7bd40001ffd3de3fa9ffffffffffffffff"),
                (x"fffffffffffffffa5287f5280fffffffffffffffffffffffff"),

                -- 3_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffff7bdea5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffdef1ce739ce7f7a94a7fffffffffffff"),
                (x"ffffffffffffffffffdef1ce739ce7f7a94a7fffffffffffff"),
                (x"ffffffffffffff4f78e718c6318c6318cfef53ffffffffffff"),
                (x"ffffffffffffe9e39c6318c6318c6318c673fa9fffffffffff"),
                (x"fffffffffffd3c718c6339cfef78e739c6319fd4ffffffffff"),
                (x"fffffffffffd3c718c6339cfef78e739c6319fd4ffffffffff"),
                (x"fffffffffffd0e339ce7f3de5295eff7bc739fd4ffffffffff"),
                (x"ffffffffffa786739cef294a3a78a51bfdef7bdea53fffffff"),
                (x"ffffffffffa787e39de57d28307a9478dfef7a9ea53fffffff"),
                (x"ffffffffffa1fc77bcaf18003078007f86f7fa9ea53fffffff"),
                (x"ffffffffffa1e9e295e318003a78007fbc31fa94a53fffffff"),
                (x"ffffffffffa1e9e295e318003a78007fbc31fa94a53fffffff"),
                (x"ffffffffffa01efa53cf1d283a7a947fbd4a3de0a53fffffff"),
                (x"ffffffffffa03de0001e78c637f9eff780007bc0a53fffffff"),
                (x"ffffffffffa529e0032005294a52940032007a94a53fffffff"),
                (x"ffffffffffa501400339c9ce739ce7ce72005014a53fffffff"),
                (x"ffffffffffa501400339c9ce739ce7ce72005014a53fffffff"),
                (x"fffffffffff8014a53339fbd4a53de9cf34a5000ffffffffff"),
                (x"ffffffffffffc1ea5333f14a529463f4f34a781fffffffffff"),
                (x"ffffffffffffc14f787428c63079ef1d1fef501fffffffffff"),
                (x"fffffffffffd3d4f79f47800307800f51fef53d4ffffffffff"),
                (x"fffffffffffd3d4f79f47800307800f51fef53d4ffffffffff"),
                (x"fffffffe94f7bdea53d47d28307a94f53d4a78e7a53fffffff"),
                (x"ffffffd0e73d3d4ef7d4a3deff7bdea529def8e7f7a9ffffff"),
                (x"fffffff86319fd4a53ddf5294a5294efa94a50e318fdffffff"),
                (x"ffffffd3bda53d4003d439ce739ce7a7a80053be39c74fffff"),
                (x"ffffffd3bda53d4003d439ce739ce7a7a80053be39c74fffff"),
                (x"ffffffd294a5294a5294f7bdef7bdef5014a7a9df78f4fffff"),
                (x"ffffffd3def501f00294a5294a5294a528319fd4a53d4fffff"),
                (x"ffffffd0e73f81f0029ea529def694a528739fd4a529ffffff"),
                (x"ffffff80e7f53ffa5294f7bc718ce7f5014a7a80ffffffffff"),
                (x"ffffff80e7f53ffa5294f7bc718ce7f5014a7a80ffffffffff"),
                (x"fffffffc00003ff003c71d294f1fdea52800001fffffffffff"),
                (x"fffffffffffffffffe9ef1ce3a0294a53fffffffffffffffff"),
                (x"fffffffffffffffffff4f7bdea0294f03fffffffffffffffff"),
                (x"ffffffffffffffffffe0a7bd40000007ffffffffffffffffff"),
                (x"ffffffffffffffffffe0a7bd40000007ffffffffffffffffff"),
                (x"ffffffffffffffffffff00c6707fffffffffffffffffffffff"),

                -- 3_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffdef7bdea5294a53fffffffffffffffff"),
                (x"ffffffffffffffef78e718c6318ce7f7a94a7fffffffffffff"),
                (x"ffffffffffffffef78e718c6318ce7f7a94a7fffffffffffff"),
                (x"fffffffffffffc718c6318c6739ce739cfef53ffffffffffff"),
                (x"ffffffffffff9e37bfc318c6319ce739ce73fa9fffffffffff"),
                (x"fffffffffffbca518c7e18c6318c6339ce739e9fffffffffff"),
                (x"fffffffffffbca518c7e18c6318c6339ce739e9fffffffffff"),
                (x"ffffffffffa1683f79e3f1cfef1c6319fc739fd4ffffffffff"),
                (x"ffffffffffa1403003cf1fbde3fbde39fdef1fd4ffffffffff"),
                (x"ffffffffffa0c0f0029ef0c63a53def1cfef7bdea53fffffff"),
                (x"ffffffffffa3c0f0029ef7bcf1be94a78fef7bdea53fffffff"),
                (x"ffffffffff03e9ea53def7bdef79ef783def7bdea53fffffff"),
                (x"ffffffffff03e9ea53def7bdef79ef783def7bdea53fffffff"),
                (x"fffffffffff83def78000529ef7bdef029ef7bdea53fffffff"),
                (x"fffffffffff800000000c8014f7bdea03def7bd4ffffffffff"),
                (x"fffffffffff80e739f39c8014a5000a7bd4a7bd4ffffffffff"),
                (x"fffffffffff80e739e73c800fa5000a53d4a7a9fffffffffff"),
                (x"fffffffffff80e739e73c800fa5000a53d4a7a9fffffffffff"),
                (x"fffffffffff8ca518e93f3dfea5000a5294a529fffffffffff"),
                (x"ffffffffffa140f7bc747fbdea5000a5294a7bffffffffffff"),
                (x"ffffffffffa0c0f001f4f7bdea5000a5294a7fffffffffffff"),
                (x"fffffffffff800fa51f4f7bd4a0294a53fffffffffffffffff"),
                (x"fffffffffff800fa51f4f7bd4a0294a53fffffffffffffffff"),
                (x"ffffffffffffc00a5294a000007694a03fffffffffffffffff"),
                (x"fffffffffffffffa5294a529eed0e7f03fffffffffffffffff"),
                (x"fffffffffffffffa53c7f77b4a78631f81ffffffffffffffff"),
                (x"fffffffffffffffa50e7a52943d3de3f81ffffffffffffffff"),
                (x"fffffffffffffffa50e7a52943d3de3f81ffffffffffffffff"),
                (x"fffffffffffffffa53d4f1cfdf1e94f501ffffffffffffffff"),
                (x"fffffffffffffffa53c718c7da7a94a028007fffffffffffff"),
                (x"fffffffffffffffffe9e19cf4efa94053c007fffffffffffff"),
                (x"fffffffffffffffffe8000014a5000a53d4a7fffffffffffff"),
                (x"fffffffffffffffffe8000014a5000a53d4a7fffffffffffff"),
                (x"fffffffffffffffffe94a0000002943fa8007fffffffffffff"),
                (x"ffffffffffffffffffc7f5280a1ce7f528007fffffffffffff"),
                (x"fffffffffffffffffe9ea529405294a529ffffffffffffffff"),
                (x"fffffffffffffffa53c7f529ff8000a7bdffffffffffffffff"),
                (x"fffffffffffffffa53c7f529ff8000a7bdffffffffffffffff"),
                (x"fffffffffffffffffffffffff053de3d29ffffffffffffffff"),

                -- 3_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffef7bdef7bdef7bfffffffffffffffff"),
                (x"ffffffffffffffff7bc739ce739ce739fdef7fffffffffffff"),
                (x"ffffffffffffffff7bc739ce739ce739fdef7fffffffffffff"),
                (x"ffffffffffffffe39ce318c6318c6319ce73fbffffffffffff"),
                (x"ffffffffffffe8718c6318c6318c6318ce739e9fffffffffff"),
                (x"fffffffffffd3c318c6318c6318c6318c6739fd4ffffffffff"),
                (x"fffffffffffd3c318c6318c6318c6318c6739fd4ffffffffff"),
                (x"fffffffffffd0e318c6318c6318c6318c6739cf4ffffffffff"),
                (x"ffffffffffa786318ce318c6318c6318ce739cfea53fffffff"),
                (x"ffffffffffa1c6318ce718c6318c6319ce739cfea53fffffff"),
                (x"ffffffffffa0ce318ce739ce739ce739ce739cfea53fffffff"),
                (x"ffffffffffa0fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa0fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa1fc318ce739ce739ce739ce739fdea53fffffff"),
                (x"ffffffffffa7bc718c7e39ce739ce73f8e739fdea53fffffff"),
                (x"ffffffffffa7bde39c7e39ce739ce7f78e73fbdea53fffffff"),
                (x"fffffffffffd3de39ce7f1ce739ce7f1ce73fbd4a53fffffff"),
                (x"fffffffffffd3de39ce7f1ce739ce7f1ce73fbd4a53fffffff"),
                (x"fffffffffffd3def78e7f7bc739fdef1cfef7bd4ffffffffff"),
                (x"ffffffffffffe9ef7bc73d29ef7a9439fdef7a9fffffffffff"),
                (x"ffffffffffffff4f7bdef5294a7a94f7bdef53ffffffffffff"),
                (x"ffffffffffffff4a529df77b4a529405294a7a9fffffffffff"),
                (x"ffffffffffffff4a529df77b4a529405294a7a9fffffffffff"),
                (x"ffffffffffffe9ef7a9df7bde1fbdef77bef1fd4ffffffffff"),
                (x"ffffffffffffe87f7a9df7bdef7bdef7a9ef78fea53fffffff"),
                (x"fffffffffffd29ef7a94efbdef53def769ef53d4a529ffffff"),
                (x"ffffffffffa53d4f7a94a529def694a529ef53dea529ffffff"),
                (x"ffffffffffa53d4f7a94a529def694a529ef53dea529ffffff"),
                (x"ffffffffffa529ef7bc0a5294a5294a53c000294a53fffffff"),
                (x"ffffffffff053b4a5280a5294ef7bda5294a53b4a53fffffff"),
                (x"fffffffffffd29def694f1cfea78e719fc005294ffffffffff"),
                (x"fffffffffff8294a5014a7bd400294f7a800001fffffffffff"),
                (x"fffffffffff8294a5014a7bd400294f7a800001fffffffffff"),
                (x"fffffffffffffe000014a5294078e73d01ffffffffffffffff"),
                (x"ffffffffffffffffffe0a5280f5294f781ffffffffffffffff"),
                (x"ffffffffffffffffffff00000f1ce7a03fffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a53de07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a53de07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0a529407ffffffffffffffffff"),

                -- 3_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294f7bdef7bfffffffffffffffff"),
                (x"ffffffffffffff4a53de38c6318c6339fdef7fffffffffffff"),
                (x"ffffffffffffff4a53de38c6318c6339fdef7fffffffffffff"),
                (x"ffffffffffffe9e39ce739ce738c6318c673fbffffffffffff"),
                (x"fffffffffffd3c739ce739ce318c631f9e31bfdfffffffffff"),
                (x"fffffffffffd0e739ce718c6318c63f0c65295ffffffffffff"),
                (x"fffffffffffd0e739ce718c6318c63f0c65295ffffffffffff"),
                (x"ffffffffffa78e7f78e319cfef1fde1bfc31d0b4ffffffffff"),
                (x"ffffffffffa78fef78e7f7bc7f78637f803180b4ffffffffff"),
                (x"fffffffe94f7bde39cfef529418fdef500f78074ffffffffff"),
                (x"fffffffe94f7bde39fd4a3de37fbdef500f781f4ffffffffff"),
                (x"fffffffe94f7bdef780f7fbdef7bdef7a9ef51e0ffffffffff"),
                (x"fffffffe94f7bdef780f7fbdef7bdef7a9ef51e0ffffffffff"),
                (x"fffffffe94f7bdea501ef7bdef5000003def781fffffffffff"),
                (x"ffffffffffa7bdef7814f7bdea0339000000001fffffffffff"),
                (x"ffffffffffa7bd4f7bd405294a0339ce4e739c1fffffffffff"),
                (x"fffffffffffd3d4f7a9405294783399cce739c1fffffffffff"),
                (x"fffffffffffd3d4f7a9405294783399cce739c1fffffffffff"),
                (x"fffffffffffd294a529405294f3fde9d0652947fffffffffff"),
                (x"fffffffffffffd4a529405294f79ef18def780b4ffffffffff"),
                (x"ffffffffffffff4a529405294f7bdef3c0f78074ffffffffff"),
                (x"fffffffffffffffffe94a0014a7bdef3e8f7801fffffffffff"),
                (x"fffffffffffffffffe94a0014a7bdef3e8f7801fffffffffff"),
                (x"fffffffffffffff00294a528000294a5280003ffffffffffff"),
                (x"fffffffffffffe0f78f4efbd4a5294a03fffffffffffffffff"),
                (x"ffffffffffffff439c7ea77beefbdef53fffffffffffffffff"),
                (x"ffffffffffffc1e39fdea529eef8e73d014a7fffffffffffff"),
                (x"ffffffffffffc1e39fdea529eef8e73d014a7fffffffffffff"),
                (x"ffffffffffffc14f78e7f5294a78e73fa9ef53ffffffffffff"),
                (x"ffffffffffffc1439fdda0000a53def529ef53ffffffffffff"),
                (x"fffffffffffffe0f7bb4a7bc7a53bded014a03ffffffffffff"),
                (x"fffffffffffffe0a5294a7bde053def501ffffffffffffffff"),
                (x"fffffffffffffe0a5294a7bde053def501ffffffffffffffff"),
                (x"fffffffffffffff00294a529405294a53fffffffffffffffff"),
                (x"fffffffffffffffa501400000a50e719ffffffffffffffffff"),
                (x"fffffffffffffffa529400014a1fdef53fffffffffffffffff"),
                (x"fffffffffffffff00000f8000a7a94a501ffffffffffffffff"),
                (x"fffffffffffffff00000f8000a7a94a501ffffffffffffffff"),
                (x"fffffffffffffffffffffffff07bde39c1ffffffffffffffff"),

                -- 3_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffff318c6a5294a7ffffffffffffffffff"),
                (x"ffffffffffffffffffdef1ce739ce731a94a7fffffffffffff"),
                (x"ffffffffffffffffffdef1ce739ce731a94a7fffffffffffff"),
                (x"ffffffffffffff4f78e718c6318c6318cfef53ffffffffffff"),
                (x"ffffffffffffe9e39c6318c6318c6318c673fa9fffffffffff"),
                (x"fffffffffffd3c718c6339cfef78e739c6319fd4ffffffffff"),
                (x"fffffffffffd3c718c6339cfef78e739c6319fd4ffffffffff"),
                (x"fffffffffffd0e339ce7f3de5295eff7bc739fd4ffffffffff"),
                (x"ffffffffffa786739cef294a3a78a51bfdef7bdea53fffffff"),
                (x"ffffffffffa787e39de57d28307a9478dfef7a9ea53fffffff"),
                (x"ffffffffffa1fc77bcaf18003078007f86f7fa9ea53fffffff"),
                (x"ffffffffffa1e9e295e318003a78007fbc31fa94a53fffffff"),
                (x"ffffffffffa1e9e295e318003a78007fbc31fa94a53fffffff"),
                (x"ffffffffffa01efa53cf1d283a7a947fbd4a3de0a53fffffff"),
                (x"ffffffffffa03de0001e78c637f9eff780007bc0a53fffffff"),
                (x"ffffffffffa529e0032005294a52940032007a94a53fffffff"),
                (x"ffffffffffa501400339c9ce739ce7ce72005014a53fffffff"),
                (x"ffffffffffa501400339c9ce739ce7ce72005014a53fffffff"),
                (x"fffffffffff8014a53339fbd4a53de9cf34a5000ffffffffff"),
                (x"ffffffffffffc1ea5333f14a529463f4f34a781fffffffffff"),
                (x"ffffffffffffc14f787428c63079ef1d1fef501fffffffffff"),
                (x"fffffffffffd3d4f79f47800307800f51fef53d4ffffffffff"),
                (x"fffffffffffd3d4f79f47800307800f51fef53d4ffffffffff"),
                (x"ffffffffffa1cfea53d47d28307a94f53d4a7bdef7bdffffff"),
                (x"fffffffe94f1fdeef694a3deff7bdea53ddefa9e39cfefffff"),
                (x"ffffffffde18cfea529eed294a5294f77d4a53c739c7ea7fff"),
                (x"ffffffd0633fbb40029ea1ce739ce73d3c0053d4a53b4a7fff"),
                (x"ffffffd0633fbb40029ea1ce739ce73d3c0053d4a53b4a7fff"),
                (x"ffffffd0e7ed29ea5014f7bdef7bdef5294a5294a5294fffff"),
                (x"fffffffe94a53c718e94a5294a5294a528007c14f7bd4fffff"),
                (x"ffffffffffa53c739e94a529def694a7a8007c1e39cf4fffff"),
                (x"fffffffffff829ea5014f1ce319fdef5294a7ff4f78e0fffff"),
                (x"fffffffffff829ea5014f1ce319fdef5294a7ff4f78e0fffff"),
                (x"ffffffffffffc0000294a7bc7f529419fc007fe00001ffffff"),
                (x"fffffffffffffffffff4a5280a0ce7f7a9ffffffffffffffff"),
                (x"ffffffffffffffffffe0f5280a7bdef53fffffffffffffffff"),
                (x"ffffffffffffffffffff00000053dea03fffffffffffffffff"),
                (x"ffffffffffffffffffff00000053dea03fffffffffffffffff"),
                (x"fffffffffffffffffffffffff01c6307ffffffffffffffffff"),

                -- 3_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffdef7bdea5294a53fffffffffffffffff"),
                (x"ffffffffffffffef78e718c6318ce7f7a94a7fffffffffffff"),
                (x"ffffffffffffffef78e718c6318ce7f7a94a7fffffffffffff"),
                (x"fffffffffffffc718c6318c6739ce739cfef53ffffffffffff"),
                (x"ffffffffffff9e37bfc318c6319ce739ce73fa9fffffffffff"),
                (x"fffffffffffbca518c7e18c6318c6339ce739e9fffffffffff"),
                (x"fffffffffffbca518c7e18c6318c6339ce739e9fffffffffff"),
                (x"ffffffffffa1683f79e3f1cfef1c6319fc739fd4ffffffffff"),
                (x"ffffffffffa1403003cf1fbde3fbde39fdef1fd4ffffffffff"),
                (x"ffffffffffa0c0f0029ef0c63a53def1cfef7bdea53fffffff"),
                (x"ffffffffffa3c0f0029ef7bcf1be94a78fef7bdea53fffffff"),
                (x"ffffffffff03e9ea53def7bdef79ef783def7bdea53fffffff"),
                (x"ffffffffff03e9ea53def7bdef79ef783def7bdea53fffffff"),
                (x"fffffffffff83def78000529ef7bdef029ef7bdea53fffffff"),
                (x"fffffffffff800000000c8014f7bdea03def7bd4ffffffffff"),
                (x"fffffffffff80e739f39c8014a5000a7bd4a7bd4ffffffffff"),
                (x"fffffffffff80e739e73c800fa5000a53d4a7a9fffffffffff"),
                (x"fffffffffff80e739e73c800fa5000a53d4a7a9fffffffffff"),
                (x"fffffffffff8ca518e93f3dfea5000a5294a529fffffffffff"),
                (x"ffffffffffa140f7bc747fbdea5000a5294a7bffffffffffff"),
                (x"ffffffffffa0c0f001f4f7bdea5000a5294a7fffffffffffff"),
                (x"fffffffffff800fa51f4f7bd4a0294a53fffffffffffffffff"),
                (x"fffffffffff800fa51f4f7bd4a0294a53fffffffffffffffff"),
                (x"ffffffffffffc00a5294a000005294a501ffffffffffffffff"),
                (x"fffffffffffffffffc14a5294a7bbda1fc007fffffffffffff"),
                (x"fffffffffffffffffe9ef7bddf7694f0cf4a7fffffffffffff"),
                (x"ffffffffffffff4002873fbddf5294f78fef03ffffffffffff"),
                (x"ffffffffffffff4002873fbddf5294f78fef03ffffffffffff"),
                (x"ffffffffffffe9ea53c73fbd4a53de39fd4a03ffffffffffff"),
                (x"ffffffffffffe9ea529ef529400294ef8f4a03ffffffffffff"),
                (x"ffffffffffffc140029ded2943fa94a77c007fffffffffffff"),
                (x"fffffffffffffff0029ef5280f7a94a528007fffffffffffff"),
                (x"fffffffffffffff0029ef5280f7a94a528007fffffffffffff"),
                (x"fffffffffffffffffe94a5280a5294a501ffffffffffffffff"),
                (x"fffffffffffffffffce33d29400000a029ffffffffffffffff"),
                (x"fffffffffffffffffe9ef1cf4a0000a529ffffffffffffffff"),
                (x"fffffffffffffff00294a7bd4003ff0001ffffffffffffffff"),
                (x"fffffffffffffff00294a7bd4003ff0001ffffffffffffffff"),
                (x"fffffffffffffff000e7f7bc0fffffffffffffffffffffffff"),

                -- 4_character_0_0
                (x"fffffffffffffffffe94a5294a5294a529ffffffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a53ffffffffffff"),
                (x"fffffffffffd28c6318c6318c6318c633cc63294ffffffffff"),
                (x"fffffffffffd28c6318c6318c6318c633cc63294ffffffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"fffffffffffd28c6318c6318c6318c6318c63294ffffffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318ca53fffffff"),
                (x"fffffffe94a328c6318c6318c6318c6318c6328ca529ffffff"),
                (x"fffffffe94a518c633cc67bcc633def3194a3194a529ffffff"),
                (x"fffffffe94a51946318c67bde6318c6318c65194a529ffffff"),
                (x"fffffffe94a52946318ca318c6318c6518c65294a529ffffff"),
                (x"fffffffe94a52946318ca318c6318c6518c65294a529ffffff"),
                (x"fffffffe94a5194a5194a318c6518c6528c65294a529ffffff"),
                (x"ffffffffff05194a5194a528ca518ca5294a5294003fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294003fffffff"),
                (x"fffffffffff8294a5194a5294a5294a5294a5280ffffffffff"),
                (x"fffffffffff8294a5194a5294a5294a5294a5280ffffffffff"),
                (x"ffffffffffffc14a5194a3194a3294a5294a501fffffffffff"),
                (x"fffffffffffffe0a528ca3194a3294a5294a03ffffffffffff"),
                (x"ffffffffffff9e400294a5294a5294a5280011feffffffffff"),
                (x"ffffffffff7902121000a5294a5294a0004204247bffffffff"),
                (x"ffffffffff7902121000a5294a5294a0004204247bffffffff"),
                (x"ffffffffff2842129463052940529400c7de8421297fffffff"),
                (x"fffffffdef094a4a53c3f0c6318c63f0fd4a10a5085fffffff"),
                (x"ffffffffde20425a53de18c6318c631fbd4a1421213dffffff"),
                (x"fffffffd8c4b19e003a318c6318c6318fa00798c4a59ffffff"),
                (x"fffffffd8c4b19e003a318c6318c6318fa00798c4a59ffffff"),
                (x"fffffffc004dd20ef7ddf7bc318fdef77dde81374a41ffffff"),
                (x"ffffffffff0000cef7bdf5294a5294f77bdeb000003fffffff"),
                (x"fffffffffffffe0ef4e718c67e9c6319cfde83ffffffffffff"),
                (x"fffffffffffffffef4e718c67e9c6319cfdeffffffffffffff"),
                (x"fffffffffffffffef4e718c67e9c6319cfdeffffffffffffff"),
                (x"fffffffffffffffef7a739cfdef4e739fbdeffffffffffffff"),
                (x"fffffffffffffff003bdef7bd077bdef7a007fffffffffffff"),
                (x"fffffffffffffff003bd3f7bd077bd3f7a007fffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc1df77a0f83bdf741ffffffffffffffff"),

                -- 4_character_0_1
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a5294ffffffffff"),
                (x"ffffffffffffe946319e6318c6318c6318c6318ca529ffffff"),
                (x"ffffffffffffe946319e6318c6318c6318c6318ca529ffffff"),
                (x"fffffffffffd28c6318c6318c632946318c63294a53fffffff"),
                (x"fffffffffffd18c6318cf318c63294a33d4a3194a53fffffff"),
                (x"ffffffffffa51946318c6528cf52944d194a518ca53fffffff"),
                (x"ffffffffffa51946318c6528cf52944d194a518ca53fffffff"),
                (x"ffffffffffa528c6318c6528c65129ba68c6528ca53fffffff"),
                (x"ffffffffffa518ca518c6528ca26f7bdee94b294a53fffffff"),
                (x"ffffffffffa3294631946528ca5ef7bdef7ba694a53fffffff"),
                (x"ffffffffffa529463294652944b18cf32f7bdc14ffffffffff"),
                (x"ffffffffff05294a5294a5294bb18ca5297bdc1fffffffffff"),
                (x"ffffffffff05294a5294a5294bb18ca5297bdc1fffffffffff"),
                (x"ffffffffff05294a5294a3189ba4a5002f7bdc1fffffffffff"),
                (x"fffffffffffd294a5289a3197ba484002f7bdc1fffffffffff"),
                (x"fffffffffff8294a5289a5297bdc84632f7bdc1fffffffffff"),
                (x"ffffffffffffc14a5294a5297bdc84632ec63194ffffffffff"),
                (x"ffffffffffffc14a5294a5297bdc84632ec63194ffffffffff"),
                (x"fffffffffffffe0a5294a2537bdd8cbdd9ef798cffffffffff"),
                (x"fffffffffffffff00294a3197bde94633cc6329fffffffffff"),
                (x"fffffffffffffffffe94a528cbde94a318c653ffffffffffff"),
                (x"ffffffffffffffffffc4214be6318ca5294a7fffffffffffff"),
                (x"ffffffffffffffffffc4214be6318ca5294a7fffffffffffff"),
                (x"ffffffffffffffff78810908fed294603dffffffffffffffff"),
                (x"ffffffffffffffe295e57bde5f0c63633bef7fffffffffffff"),
                (x"ffffffffffffffe7bc81094aff786365bdef7fffffffffffff"),
                (x"ffffffffffffffe210bef318c003deeb19ef7fffffffffffff"),
                (x"ffffffffffffffe210bef318c003deeb19ef7fffffffffffff"),
                (x"fffffffffffffe029597ba537ba4001d99ef7fffffffffffff"),
                (x"fffffffffffffe0632f7bdef7bdc00f599ef7fffffffffffff"),
                (x"fffffffffffffff00137ba537ba400edbdffffffffffffffff"),
                (x"fffffffffffffffffc006318c000e73f7fffffffffffffffff"),
                (x"fffffffffffffffffc006318c000e73f7fffffffffffffffff"),
                (x"fffffffffffffffffc1def7bde9ce7ef7fffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7bd38ce7efffffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7a719fbdffffffffffffffffffff"),
                (x"ffffffffffffffffffff077a318c00ffffffffffffffffffff"),
                (x"ffffffffffffffffffff077a318c00ffffffffffffffffffff"),
                (x"ffffffffffffffffffff077be2f800ffffffffffffffffffff"),

                -- 4_character_0_2
                (x"fffffffffffffffffe94a5294a5294a529ffffffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c65294a53ffffffffffff"),
                (x"fffffffffffd28c633cc6318c6318c6318c65294ffffffffff"),
                (x"fffffffffffd28c633cc6318c6318c6318c65294ffffffffff"),
                (x"ffffffffffa518c6319e6528c6318c6319ef3194a53fffffff"),
                (x"fffffffffffd28c6318ca528cf329467a8c63294ffffffffff"),
                (x"ffffffffffa518ca5194a529465294a3194a3194a53fffffff"),
                (x"ffffffffffa518ca5194a529465294a3194a3194a53fffffff"),
                (x"ffffffffffa318ca519462534a518c4d194a328ca53fffffff"),
                (x"fffffffe94a328ca528cbdee9a32f7ba694a52946329ffffff"),
                (x"fffffffe94651944a697bdef765ef7bde894d294a529ffffff"),
                (x"fffffffe94a5194bdd37bdef7bdef7bdd37bd194a529ffffff"),
                (x"fffffffe94a52946319e65ef7bdef76798c65294a529ffffff"),
                (x"fffffffe94a52946319e65ef7bdef76798c65294a529ffffff"),
                (x"fffffffe94a528c63194a5297bde94a518c63294a529ffffff"),
                (x"ffffffffff0268cbdca005ef7bdef7000b7bb289003fffffff"),
                (x"ffffffffff0268cbdc8005ef7bdef700097bb289003fffffff"),
                (x"fffffffffff8294bdc8c65ef7bdef763097bd280ffffffffff"),
                (x"fffffffffff8294bdc8c65ef7bdef763097bd280ffffffffff"),
                (x"ffffffffffffc14bdc8c6318cbb18c63097bd01fffffffffff"),
                (x"fffffffffffbca0632f767bdea7bde65eec600afffffffffff"),
                (x"ffffffffff79025a518cf318ca318cf3194a14247bffffffff"),
                (x"fffffffdef28424a528c63194bd18c63294a1021295fffffff"),
                (x"fffffffdef28424a528c63194bd18c63294a1021295fffffff"),
                (x"ffffffbc84215e429694a528c63294a5285291e52108ffffff"),
                (x"fffff797def10af297be18c7ef78631fba52bca4f7bc57ffff"),
                (x"fffff7b1294b09e003d41d28cb32941d3c00788c4a52c7ffff"),
                (x"fffff626f7ba580003c3a77a3677bda0fc000189bdee967fff"),
                (x"fffff626f7ba580003c3a77a3677bda0fc000189bdee967fff"),
                (x"fffff626f74deec0028318c6cb306318e80032f74a6e967fff"),
                (x"ffffff81294deecef7d4f7bccb33def53ddeb2f74a520fffff"),
                (x"fffffffc004dee0ef4fef7bde67bdef78fde82f74a41ffffff"),
                (x"ffffffffff0001fef4e718c6318c6319cfdefc00003fffffff"),
                (x"ffffffffff0001fef4e718c6318c6319cfdefc00003fffffff"),
                (x"fffffffffffffffef7a719cfdef4e719fbdeffffffffffffff"),
                (x"fffffffffffffff003a739cfd074e739fa007fffffffffffff"),
                (x"fffffffffffffff003a319cfd074e718fa007fffffffffffff"),
                (x"fffffffffffffffffc1def7a0f83bdef41ffffffffffffffff"),
                (x"fffffffffffffffffc1def7a0f83bdef41ffffffffffffffff"),
                (x"ffffffffffffffffffbdf77a0f83bdf77bffffffffffffffff"),

                -- 4_character_0_3
                (x"ffffffffffffff4a52946318c65294a53fffffffffffffffff"),
                (x"ffffffffffa52946318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf3194a53ffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf3194a53ffffffffffff"),
                (x"fffffffe94a518c6318ca318c6318c6318c6529fffffffffff"),
                (x"fffffffe94a3194f7994a318c633de6318c6329fffffffffff"),
                (x"fffffffe946329463289a529e6518c63194a3294ffffffffff"),
                (x"fffffffe946329463289a529e6518c63194a3294ffffffffff"),
                (x"fffffffe946528ca51374d28c6518c6318c65294ffffffffff"),
                (x"fffffffe94a5189bdef7ba5346518c6328c63294ffffffffff"),
                (x"fffffffe94a5137bdef7bdef46518ca3194a5194ffffffffff"),
                (x"ffffffffffa02f7bdd9e63189a518ca5194a5294ffffffffff"),
                (x"fffffffffff82f7a529463197a5294a5294a5280ffffffffff"),
                (x"fffffffffff82f7a529463197a5294a5294a5280ffffffffff"),
                (x"fffffffffff82f7bdc002a5374b294a5294a5280ffffffffff"),
                (x"fffffffffff82f7bdc0022537bb2944d294a501fffffffffff"),
                (x"fffffffffff82f7bdd8c25ef7bd2944d294a501fffffffffff"),
                (x"ffffffffffa318cbdd8c25ef7bd294a5294a03ffffffffffff"),
                (x"ffffffffffa318cbdd8c25ef7bd294a5294a03ffffffffffff"),
                (x"ffffffffff633de632f765ef7ba694a528007fffffffffffff"),
                (x"ffffffffff6518cf798ca5ef7bb294a501ffffffffffffffff"),
                (x"fffffffffffd28c63194a5ef765294a53fffffffffffffffff"),
                (x"ffffffffffffff4a52946318cf148427bfffffffffffffffff"),
                (x"ffffffffffffff4a52946318cf148427bfffffffffffffffff"),
                (x"ffffffffffffffff780ca529d79021093dffffffffffffffff"),
                (x"ffffffffffffffeef58c18c7e2bdef2bcbef7fffffffffffff"),
                (x"ffffffffffffffef7acc1fbde79421091fef7fffffffffffff"),
                (x"ffffffffffffffe6319df0000633def149ef7fffffffffffff"),
                (x"ffffffffffffffe6319df0000633def149ef7fffffffffffff"),
                (x"ffffffffffffffe632c302537ba6f7bb0a007fffffffffffff"),
                (x"ffffffffffffffe632de05ef7bdef7bdd8007fffffffffffff"),
                (x"ffffffffffffffff7add02537ba6f7ba41ffffffffffffffff"),
                (x"ffffffffffffffffffa7380006318c003fffffffffffffffff"),
                (x"ffffffffffffffffffa7380006318c003fffffffffffffffff"),
                (x"ffffffffffffffffffbd39cfdef7bde83fffffffffffffffff"),
                (x"fffffffffffffffffffd38c67ef7bd07ffffffffffffffffff"),
                (x"ffffffffffffffffffffe9ce33f7bd07ffffffffffffffffff"),
                (x"ffffffffffffffffffff00c631f400ffffffffffffffffffff"),
                (x"ffffffffffffffffffff00c631f400ffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc5f7400ffffffffffffffffffff"),

                -- 4_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a529ffffffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a53ffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a53ffffffffffff"),
                (x"fffffffffffd28c6318c6318c6318c633cc63294ffffffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"fffffffffffd28c6318c6318c6318c6318c63294ffffffffff"),
                (x"fffffffffffd28c6318c6318c6318c6318c63294ffffffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318ca53fffffff"),
                (x"fffffffe94a328c6318c6318c6318c6318c6328ca529ffffff"),
                (x"fffffffe94a518c633cc67bcc633def3194a3194a529ffffff"),
                (x"fffffffe94a51946318c67bde6318c6318c65194a529ffffff"),
                (x"fffffffe94a51946318c67bde6318c6318c65194a529ffffff"),
                (x"fffffffe94a52946318ca318c6318c6518c65294a529ffffff"),
                (x"fffffffe94a5194a5194a318c6518c6528c65294a529ffffff"),
                (x"ffffffffff05194a5194a528ca518ca5294a5294003fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294003fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294003fffffff"),
                (x"fffffffffff8294a5194a5294a5294a5294a5280ffffffffff"),
                (x"ffffffffffffc14a5194a3194a3294a5294a501fffffffffff"),
                (x"fffffffffffffc0a528ca3194a3294a5294a03ffffffffffff"),
                (x"ffffffffffff8a400294a5294a5294a5280013dfffffffffff"),
                (x"ffffffffffff8a400294a5294a5294a5280013dfffffffffff"),
                (x"fffffffffff1484ef400a5294a5294a00010849effffffffff"),
                (x"fffffffffff10a5a5063052940529407ba10843effffffffff"),
                (x"fffffffffff1484f787e18c631f8631fba108485f7bfffffff"),
                (x"ffffffffff67bdea53c318c631fbbd1fa8529484f7bfffffff"),
                (x"ffffffffff67bdea53c318c631fbbd1fa8529484f7bfffffff"),
                (x"ffffffffff03180a53be18c6318fdeef6810843e633fffffff"),
                (x"fffffffffff8000f7a9defbdeef7def781ef7bc9633fffffff"),
                (x"fffffffffffffffef7bd39cfdef7bdef7ac62520ffffffffff"),
                (x"fffffffffffffffef7bd38c63ef4e73f7bde801fffffffffff"),
                (x"fffffffffffffffef7bd38c63ef4e73f7bde801fffffffffff"),
                (x"fffffffffffffffef7bde9ce7ef7bdef40007fffffffffffff"),
                (x"fffffffffffffffffc1def7bd383bde83fffffffffffffffff"),
                (x"ffffffffffffffffffe0e9ce7e800007ffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc3f03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc3f03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bdde83ffffffffffffffffffffff"),

                -- 4_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a5294ffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a5294ffffffffff"),
                (x"ffffffffffffe946319e6318c6318c6318c6318ca529ffffff"),
                (x"fffffffffffd28c6318c6318c632946318c63294a53fffffff"),
                (x"fffffffffffd18c6318cf318c63294a33d4a3194a53fffffff"),
                (x"fffffffffffd18c6318cf318c63294a33d4a3194a53fffffff"),
                (x"ffffffffffa51946318c6528cf52944d194a518ca53fffffff"),
                (x"ffffffffffa528c6318c6528c65129ba68c6528ca53fffffff"),
                (x"ffffffffffa518ca518c6528ca26f7bdee94b294a53fffffff"),
                (x"ffffffffffa3294631946528ca5ef7bdef7ba694a53fffffff"),
                (x"ffffffffffa529463294652944b18cf32f7bdc14ffffffffff"),
                (x"ffffffffffa529463294652944b18cf32f7bdc14ffffffffff"),
                (x"ffffffffff05294a5294a5294bb18ca5297bdc1fffffffffff"),
                (x"ffffffffff05294a5294a3189ba4a5002f7bdc1fffffffffff"),
                (x"fffffffffffd294a5289a3197ba484002f7bdc1fffffffffff"),
                (x"fffffffffff8294a5289a5297bdc84632f7bdc1fffffffffff"),
                (x"fffffffffff8294a5289a5297bdc84632f7bdc1fffffffffff"),
                (x"ffffffffffffc14a5294a5297bdc84632ec63194ffffffffff"),
                (x"fffffffffffffe0a5294a2537bdd8cbdd9ef798cffffffffff"),
                (x"fffffffffffffff00294a3197bde94633cc6328cffffffffff"),
                (x"fffffffffffffffffe94a528cbde94a318c6529fffffffffff"),
                (x"fffffffffffffffffe94a528cbde94a318c6529fffffffffff"),
                (x"fffffffffffffff003c5214af6318ca5294a7fffffffffffff"),
                (x"fffffffffffffff000a408425f5294a03dffffffffffffffff"),
                (x"fffffffffffffe0f7884294a4a7bdef798007fffffffffffff"),
                (x"fffffffffffffe0f78af08421f77def798007fffffffffffff"),
                (x"fffffffffffffe0f78af08421f77def798007fffffffffffff"),
                (x"fffffffffffffe0a51e42bdfef0000053ac67fffffffffffff"),
                (x"fffffffffffffe0a53c5f318965ef7b83ac67fffffffffffff"),
                (x"fffffffffffffe0f7a804def74def7b828c67fffffffffffff"),
                (x"ffffffffffffffd003de025374a6f76741ffffffffffffffff"),
                (x"ffffffffffffffd003de025374a6f76741ffffffffffffffff"),
                (x"ffffffffffffffdef4e7e800c60000077fffffffffffffffff"),
                (x"fffffffffffffe0ef4e33f7bd077bdefffffffffffffffffff"),
                (x"fffffffffffffe0ef7a7ef7bd074e73f7fffffffffffffffff"),
                (x"fffffffffffffff000e33f7a0003bdf7bfffffffffffffffff"),
                (x"fffffffffffffff000e33f7a0003bdf7bfffffffffffffffff"),
                (x"fffffffffffffff003be2fbc0fffffffffffffffffffffffff"),

                -- 4_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a529ffffffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c65294a53ffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c65294a53ffffffffffff"),
                (x"fffffffffffd28c633cc6318c6318c6318c65294ffffffffff"),
                (x"ffffffffffa518c6319e6528c6318c6319ef3194a53fffffff"),
                (x"fffffffffffd28c6318ca528cf329467a8c63294ffffffffff"),
                (x"fffffffffffd28c6318ca528cf329467a8c63294ffffffffff"),
                (x"ffffffffffa518ca5194a529465294a3194a3194a53fffffff"),
                (x"ffffffffffa318ca519462534a518c4d194a328ca53fffffff"),
                (x"fffffffe94a328ca528cbdee9a32f7ba694a52946329ffffff"),
                (x"fffffffe94651944a697bdef765ef7bde894d294a529ffffff"),
                (x"fffffffe94a5194bdd37bdef7bdef7bdd37bd194a529ffffff"),
                (x"fffffffe94a5194bdd37bdef7bdef7bdd37bd194a529ffffff"),
                (x"fffffffe94a52946319e65ef7bdef76798c65294a529ffffff"),
                (x"fffffffe94a528c63194a5297bde94a518c63294a529ffffff"),
                (x"ffffffffff0268cbdca005ef7bdef7000b7bb289003fffffff"),
                (x"ffffffffff0268cbdc8005ef7bdef700097bb289003fffffff"),
                (x"ffffffffff0268cbdc8005ef7bdef700097bb289003fffffff"),
                (x"fffffffffff8294bdc8c65ef7bdef763097bd280ffffffffff"),
                (x"ffffffffffffc14bdc8c6318cbb18c63097bd01fffffffffff"),
                (x"ffffffffffff9e0632f767bdea7bde65eec603deffffffffff"),
                (x"ffffffffff79485a518cf318ca318cf3194a1424f7bfffffff"),
                (x"ffffffffff79485a518cf318ca318cf3194a1424f7bfffffff"),
                (x"fffffffdef29084a528c63194bd18c63294a0484297dffffff"),
                (x"fffffff88423ca421294a528c63294a529debc21210befffff"),
                (x"fffffff9ef291efef69e18c7ef78631fa94a11ef7bcbefffff"),
                (x"ffffffb12963ca0a53d41d28cb32941d3d4a0129633dffffff"),
                (x"ffffffb12963ca0a53d41d28cb32941d3d4a0129633dffffff"),
                (x"ffffffb1294b180a53c3a77a3677bda0c00032f74a59ffffff"),
                (x"ffffffb2f7ba41fa53a318c6cb30631f597bdee94a59ffffff"),
                (x"ffffffb129bb01fef7deefbccb33bdf7997bdd2c6301ffffff"),
                (x"ffffff81294b3ffef4e718c6361ce73f4094dd80003fffffff"),
                (x"ffffff81294b3ffef4e718c6361ce73f4094dd80003fffffff"),
                (x"fffffffc00003ffef7a718c67ef7bdef7a00001fffffffffff"),
                (x"ffffffffffffffffffa738c67383bdef7bffffffffffffffff"),
                (x"fffffffffffffffffffd18c63383bdef7fffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7bde800007ffffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7bde800007ffffffffffffffffff"),
                (x"ffffffffffffffffffffef7beeffffffffffffffffffffffff"),

                -- 4_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffff4a52946318c65294a53fffffffffffffffff"),
                (x"ffffffffffa52946318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffffffa52946318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf3194a53ffffffffffff"),
                (x"fffffffe94a518c6318ca318c6318c6318c6529fffffffffff"),
                (x"fffffffe94a3194f7994a318c633de6318c6329fffffffffff"),
                (x"fffffffe94a3194f7994a318c633de6318c6329fffffffffff"),
                (x"fffffffe946329463289a529e6518c63194a3294ffffffffff"),
                (x"fffffffe946528ca51374d28c6518c6318c65294ffffffffff"),
                (x"fffffffe94a5189bdef7ba5346518c6328c63294ffffffffff"),
                (x"fffffffe94a5137bdef7bdef46518ca3194a5194ffffffffff"),
                (x"ffffffffffa02f7bdd9e63189a518ca5194a5294ffffffffff"),
                (x"ffffffffffa02f7bdd9e63189a518ca5194a5294ffffffffff"),
                (x"fffffffffff82f7a529463197a5294a5294a5280ffffffffff"),
                (x"fffffffffff82f7bdc002a5374b294a5294a5280ffffffffff"),
                (x"fffffffffff82f7bdc0022537bb2944d294a501fffffffffff"),
                (x"fffffffffff82f7bdd8c25ef7bd2944d294a501fffffffffff"),
                (x"fffffffffff82f7bdd8c25ef7bd2944d294a501fffffffffff"),
                (x"ffffffffffa318cbdd8c25ef7bd294a5294a03ffffffffffff"),
                (x"ffffffffff633de632f765ef7ba694a528007fffffffffffff"),
                (x"ffffffffff6518cf798ca5ef7bb294a501ffffffffffffffff"),
                (x"fffffffffffd28c63194a5ef765294a53fffffffffffffffff"),
                (x"fffffffffffd28c63194a5ef765294a53fffffffffffffffff"),
                (x"ffffffffffffff4a52946318c794842f81ffffffffffffffff"),
                (x"ffffffffffffffff7814a529e284212141ffffffffffffffff"),
                (x"fffffffffffffe0633def7bd4214a5213c007fffffffffffff"),
                (x"fffffffffffffe0633def77be08421797c007fffffffffffff"),
                (x"fffffffffffffe0633def77be08421797c007fffffffffffff"),
                (x"fffffffffffffecef6800001ef3ca523e8007fffffffffffff"),
                (x"fffffffffffffecef417bdeec4b3de2fa8007fffffffffffff"),
                (x"fffffffffffffeca5017bdee9bdd2903fc007fffffffffffff"),
                (x"fffffffffffffff003acba529ba400f781deffffffffffffff"),
                (x"fffffffffffffff003acba529ba400f781deffffffffffffff"),
                (x"ffffffffffffffffffa00000c603bd39fbdeffffffffffffff"),
                (x"fffffffffffffffffffdef7a0ef4e719fa007fffffffffffff"),
                (x"ffffffffffffffffffa73f7a0ef7bd3f7a007fffffffffffff"),
                (x"ffffffffffffffffffdee8000074e719c1ffffffffffffffff"),
                (x"ffffffffffffffffffdee8000074e719c1ffffffffffffffff"),
                (x"fffffffffffffffffffffffff078a5f741ffffffffffffffff"),

                -- 4_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a529ffffffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a53ffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a53ffffffffffff"),
                (x"fffffffffffd28c6318c6318c6318c633cc63294ffffffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"fffffffffffd28c6318c6318c6318c6318c63294ffffffffff"),
                (x"fffffffffffd28c6318c6318c6318c6318c63294ffffffffff"),
                (x"ffffffffffa518c6318c6318c6318c6318c63194a53fffffff"),
                (x"ffffffffffa318c6318c6318c6318c6318c6318ca53fffffff"),
                (x"fffffffe94a328c6318c6318c6318c6318c6328ca529ffffff"),
                (x"fffffffe94a518c633cc67bcc633def3194a3194a529ffffff"),
                (x"fffffffe94a51946318c67bde6318c6318c65194a529ffffff"),
                (x"fffffffe94a51946318c67bde6318c6318c65194a529ffffff"),
                (x"fffffffe94a52946318ca318c6318c6518c65294a529ffffff"),
                (x"fffffffe94a5194a5194a318c6518c6528c65294a529ffffff"),
                (x"ffffffffff05194a5194a528ca518ca5294a5294003fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294003fffffff"),
                (x"ffffffffff05294a5294a5294a5294a5294a5294003fffffff"),
                (x"fffffffffff8294a5194a5294a5294a5294a5280ffffffffff"),
                (x"ffffffffffffc14a5194a3194a3294a5294a501fffffffffff"),
                (x"fffffffffffffe0a528ca3194a3294a5294a03dfffffffffff"),
                (x"fffffffffffffc400294a5294a5294a5280013beffffffffff"),
                (x"fffffffffffffc400294a5294a5294a5280013beffffffffff"),
                (x"ffffffffffff88108400a5294a5294a001de909df7bfffffff"),
                (x"ffffffffffff821087be052940529400c74a14a4f7bfffffff"),
                (x"fffffffffff1481087be18c7e18c631f87ef1085f7bfffffff"),
                (x"fffffffffff10852969e1f7be18c6318fd4a7bde633fffffff"),
                (x"fffffffffff10852969e1f7be18c6318fd4a7bde633fffffff"),
                (x"ffffffffff678210869defbc318c631fbb4a018c003fffffff"),
                (x"ffffffffff627def781ef7bddefbdeef69ef0000ffffffffff"),
                (x"fffffffffff8129633bdef7bdef4e73f7bdeffffffffffffff"),
                (x"ffffffffffffc00ef7bd39cfde8c633f7bdeffffffffffffff"),
                (x"ffffffffffffc00ef7bd39cfde8c633f7bdeffffffffffffff"),
                (x"fffffffffffffff0001def7bde9ce7ef7bdeffffffffffffff"),
                (x"ffffffffffffffffffe0ef7a03f7bdef41ffffffffffffffff"),
                (x"ffffffffffffffffffff00000e9ce7e83fffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f0fde07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f0fde07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0ef7de07ffffffffffffffffff"),

                -- 4_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a528c6318ca5294a7fffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a5294ffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c63194a5294ffffffffff"),
                (x"ffffffffffffe946319e6318c6318c6318c6318ca529ffffff"),
                (x"fffffffffffd28c6318c6318c632946318c63294a53fffffff"),
                (x"fffffffffffd18c6318cf318c63294a33d4a3194a53fffffff"),
                (x"fffffffffffd18c6318cf318c63294a33d4a3194a53fffffff"),
                (x"ffffffffffa51946318c6528cf52944d194a518ca53fffffff"),
                (x"ffffffffffa528c6318c6528c65129ba68c6528ca53fffffff"),
                (x"ffffffffffa518ca518c6528ca26f7bdee94b294a53fffffff"),
                (x"ffffffffffa3294631946528ca5ef7bdef7ba694a53fffffff"),
                (x"ffffffffffa529463294652944b18cf32f7bdc14ffffffffff"),
                (x"ffffffffffa529463294652944b18cf32f7bdc14ffffffffff"),
                (x"ffffffffff05294a5294a5294bb18ca5297bdc1fffffffffff"),
                (x"ffffffffff05294a5294a3189ba4a5002f7bdc1fffffffffff"),
                (x"fffffffffffd294a5289a3197ba484002f7bdc1fffffffffff"),
                (x"fffffffffff8294a5289a5297bdc84632f7bdc1fffffffffff"),
                (x"fffffffffff8294a5289a5297bdc84632f7bdc1fffffffffff"),
                (x"ffffffffffffc14a5294a5297bdc84632ec63194ffffffffff"),
                (x"fffffffffffffe0a5294a2537bdd8cbdd9ef798cffffffffff"),
                (x"fffffffffffffff00294a3197bde94633cc6328cffffffffff"),
                (x"fffffffffffffffffe94a528cbde94a318c6529fffffffffff"),
                (x"fffffffffffffffffe94a528cbde94a318c6529fffffffffff"),
                (x"fffffffffffffff000a42fbde6318ca5294a7fffffffffffff"),
                (x"fffffffffffffe02942123dfdf5294483dffffffffffffffff"),
                (x"ffffffffffffffe7bc840f7be18fde67bbef7fffffffffffff"),
                (x"ffffffffffffc0f210212f7bda0d8cb7bac67fffffffffffff"),
                (x"ffffffffffffc0f210212f7bda0d8cb7bac67fffffffffffff"),
                (x"ffffffffffffc05f79ef27bd4f798c677c94b3ffffffffffff"),
                (x"ffffffffffffc1e4a6f748000f798cb77c9483ffffffffffff"),
                (x"fffffffffffffe04a6f7bdee9f758cb780007fffffffffffff"),
                (x"fffffffffffffe063137bdef701d8cb741ffffffffffffffff"),
                (x"fffffffffffffe063137bdef701d8cb741ffffffffffffffff"),
                (x"fffffffffffffff0000c4dee900c63677fffffffffffffffff"),
                (x"fffffffffffffff003bd00000e9fbdef7fffffffffffffffff"),
                (x"fffffffffffffffef7bd00000e9c6319ffffffffffffffffff"),
                (x"fffffffffffffff0001de8000074e7ef41ffffffffffffffff"),
                (x"fffffffffffffff0001de8000074e7ef41ffffffffffffffff"),
                (x"fffffffffffffffffffffffff077de2f81ffffffffffffffff"),

                -- 4_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94a5294a5294a529ffffffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c65294a53ffffffffffff"),
                (x"ffffffffffffff4a528c6318c6318c65294a53ffffffffffff"),
                (x"fffffffffffd28c633cc6318c6318c6318c65294ffffffffff"),
                (x"ffffffffffa518c6319e6528c6318c6319ef3194a53fffffff"),
                (x"fffffffffffd28c6318ca528cf329467a8c63294ffffffffff"),
                (x"fffffffffffd28c6318ca528cf329467a8c63294ffffffffff"),
                (x"ffffffffffa518ca5194a529465294a3194a3194a53fffffff"),
                (x"ffffffffffa318ca519462534a518c4d194a328ca53fffffff"),
                (x"fffffffe94a328ca528cbdee9a32f7ba694a52946329ffffff"),
                (x"fffffffe94651944a697bdef765ef7bde894d294a529ffffff"),
                (x"fffffffe94a5194bdd37bdef7bdef7bdd37bd194a529ffffff"),
                (x"fffffffe94a5194bdd37bdef7bdef7bdd37bd194a529ffffff"),
                (x"fffffffe94a52946319e65ef7bdef76798c65294a529ffffff"),
                (x"fffffffe94a528c63194a5297bde94a518c63294a529ffffff"),
                (x"ffffffffff0268cbdca005ef7bdef7000b7bb289003fffffff"),
                (x"ffffffffff0268cbdc8005ef7bdef700097bb289003fffffff"),
                (x"ffffffffff0268cbdc8005ef7bdef700097bb289003fffffff"),
                (x"fffffffffff8294bdc8c65ef7bdef763097bd280ffffffffff"),
                (x"ffffffffffffc14bdc8c6318cbb18c63097bd01fffffffffff"),
                (x"ffffffffffffbc0632f767bdea7bde65eec601feffffffffff"),
                (x"fffffffffff1025a518cf318ca318cf3194a14857bffffffff"),
                (x"fffffffffff1025a518cf318ca318cf3194a14857bffffffff"),
                (x"ffffffffde29081a528c63194bd18c63294a1084295fffffff"),
                (x"fffffff8a52042f29694a528c63294a529ef10af2109efffff"),
                (x"fffffff8a57bde4a529e18c7ef78631fa9ded1e4295fefffff"),
                (x"ffffffffde62520a53d41d28cb32941d3d4a00af6312cfffff"),
                (x"ffffffffde62520a53d41d28cb32941d3d4a00af6312cfffff"),
                (x"fffffffd8c4deec00003a77a3677bda0fd4a018c4a52cfffff"),
                (x"fffffffd8c4a6f7bdd9d18c6cb306318fb4a7c09bdeecfffff"),
                (x"fffffffc0063137bdd9ef77acb33deefbddefc0cbdd2cfffff"),
                (x"ffffffffff001974a41d39ce361c6319cfdeffec4a520fffff"),
                (x"ffffffffff001974a41d39ce361c6319cfdeffec4a520fffff"),
                (x"ffffffffffffc00003bdef7bde9c6319fbdeffe00001ffffff"),
                (x"ffffffffffffffffffbdef7a039c6339fbffffffffffffffff"),
                (x"fffffffffffffffffffdef7a038c631f7fffffffffffffffff"),
                (x"ffffffffffffffffffff00000ef7bde83fffffffffffffffff"),
                (x"ffffffffffffffffffff00000ef7bde83fffffffffffffffff"),
                (x"fffffffffffffffffffffffffefbbdefffffffffffffffffff"),

                -- 4_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffff4a52946318c65294a53fffffffffffffffff"),
                (x"ffffffffffa52946318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffffffa52946318c6318c6318c65294a7fffffffffffff"),
                (x"ffffffd2946318c6318c6318c6318cf3194a53ffffffffffff"),
                (x"fffffffe94a518c6318ca318c6318c6318c6529fffffffffff"),
                (x"fffffffe94a3194f7994a318c633de6318c6329fffffffffff"),
                (x"fffffffe94a3194f7994a318c633de6318c6329fffffffffff"),
                (x"fffffffe946329463289a529e6518c63194a3294ffffffffff"),
                (x"fffffffe946528ca51374d28c6518c6318c65294ffffffffff"),
                (x"fffffffe94a5189bdef7ba5346518c6328c63294ffffffffff"),
                (x"fffffffe94a5137bdef7bdef46518ca3194a5194ffffffffff"),
                (x"ffffffffffa02f7bdd9e63189a518ca5194a5294ffffffffff"),
                (x"ffffffffffa02f7bdd9e63189a518ca5194a5294ffffffffff"),
                (x"fffffffffff82f7a529463197a5294a5294a5280ffffffffff"),
                (x"fffffffffff82f7bdc002a5374b294a5294a5280ffffffffff"),
                (x"fffffffffff82f7bdc0022537bb2944d294a501fffffffffff"),
                (x"fffffffffff82f7bdd8c25ef7bd2944d294a501fffffffffff"),
                (x"fffffffffff82f7bdd8c25ef7bd2944d294a501fffffffffff"),
                (x"ffffffffffa318cbdd8c25ef7bd294a5294a03ffffffffffff"),
                (x"ffffffffff633de632f765ef7ba694a528007fffffffffffff"),
                (x"ffffffffff6518cf798ca5ef7bb294a501ffffffffffffffff"),
                (x"fffffffffffd28c63194a5ef765294a53fffffffffffffffff"),
                (x"fffffffffffd28c63194a5ef765294a53fffffffffffffffff"),
                (x"ffffffffffffff4a52946318cf78a52141ffffffffffffffff"),
                (x"ffffffffffffffff7809a529eed084084a007fffffffffffff"),
                (x"ffffffffffffffeef7ccf0c63f1421211fef7fffffffffffff"),
                (x"fffffffffffffecef7d660c74e94a50848f783ffffffffffff"),
                (x"fffffffffffffecef7d660c74e94a50848f783ffffffffffff"),
                (x"ffffffffffffd89f7bac67bdea78847bfc5283ffffffffffff"),
                (x"ffffffffffffc09f7bb667bde00129bdd3ef03ffffffffffff"),
                (x"fffffffffffffe0003d6677be4def7bdd2007fffffffffffff"),
                (x"fffffffffffffff003b661ce0bdef7ba58007fffffffffffff"),
                (x"fffffffffffffff003b661ce0bdef7ba58007fffffffffffff"),
                (x"ffffffffffffffffffac18c604dd296001ffffffffffffffff"),
                (x"ffffffffffffffffffbde9cfd00000ef41ffffffffffffffff"),
                (x"fffffffffffffffffce319cfd00000ef7bffffffffffffffff"),
                (x"fffffffffffffff003bd3f7a0003bde801ffffffffffffffff"),
                (x"fffffffffffffff003bd3f7a0003bde801ffffffffffffffff"),
                (x"fffffffffffffff003c5f77a0fffffffffffffffffffffffff"),

                -- 5_character_0_0
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffe9def5ce739ce739ce739ddef69fffffffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b9ae739dda53fffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b9ae739dda53fffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad6b5cd6b9ceef69ffffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae739ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ae735ce739d4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4fffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae735cd73bb4fffff"),
                (x"ffffffd3bdeb9cd6b5ad6b5ad6b5ad6b5ad6b9aeef7b4fffff"),
                (x"ffffffd294ef7ae739cd6b5ad6b5ad6b5ae73bbdef694fffff"),
                (x"ffffffd294ef7ae739cd6b5ad6b5ad6b5ae73bbdef694fffff"),
                (x"fffffffe94ef7bdef7ae739ce739ce73bbdef7bdef69ffffff"),
                (x"ffffffffffa53bdef7bdef7bdef7bdef7bdef7bda53bffffff"),
                (x"ffffffffffef694a53bdef7bdef7bdef7b4a529dffffffffff"),
                (x"ffffffffffff7b4a5294a77bdef7bda5294a5280ffffffffff"),
                (x"ffffffffffff7b4a5294a77bdef7bda5294a5280ffffffffff"),
                (x"ffffffffffffc14ef7b4ef7bdef7bded3bded01fffffffffff"),
                (x"fffffffffffffe0a53bdef7bdef7bded294a03ffffffffffff"),
                (x"ffffffffffffe94a529da77b4ed3bda5294a529fffffffffff"),
                (x"fffffffffffd3b4ef7b4a5294a5294a53bded3b4ffffffffff"),
                (x"fffffffffffd3b4ef7b4a5294a5294a53bded3b4ffffffffff"),
                (x"ffffffffffa77ddef7dee8014a5000efbddef7dda53fffffff"),
                (x"ffffffffff07bdea53def7bdef7bdef7bd4a7bde003fffffff"),
                (x"fffffffd8c4829da53bef7bd30cfdef7bb4a76804a59ffffff"),
                (x"fffffffd8c4dc00a53bef7bdef7bdef7bb4a00174a59ffffff"),
                (x"fffffffd8c4dc00a53bef7bdef7bdef7bb4a00174a59ffffff"),
                (x"fffffffc004dd20a529defbc1987deef694a01374a41ffffff"),
                (x"ffffffffff00014a53b4a529da7694a53b4a5000003fffffff"),
                (x"ffffffffffffff4a53bef7bdef7bdef7bb4a53ffffffffffff"),
                (x"fffffffffffffffa529df7bdef7bdef7694a7fffffffffffff"),
                (x"fffffffffffffffa529df7bdef7bdef7694a7fffffffffffff"),
                (x"fffffffffffffffe73bdef7bde77bdef7bce7fffffffffffff"),
                (x"fffffffffffffff003ae739dd075ce73ba007fffffffffffff"),
                (x"fffffffffffffff0038e777bc073bd73b8007fffffffffffff"),
                (x"fffffffffffffffffc1cef7a0f83bdef01ffffffffffffffff"),
                (x"fffffffffffffffffc1cef7a0f83bdef01ffffffffffffffff"),
                (x"fffffffffffffffffc0000000f80000001ffffffffffffffff"),

                -- 5_character_0_1
                (x"fffffffffffffffffffffd294ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffe94ef7ae735ad6b5ae73bb4ffffffffff"),
                (x"ffffffffffffff4ef7ae6b5ad6b5ad6b5ad6b5dda53fffffff"),
                (x"ffffffffffffff4ef7ae6b5ad6b5ad6b5ad6b5dda53fffffff"),
                (x"fffffffffffd3bd739ad6b5ad6b5ad6b5ad6b5aea53fffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b5ae777b4a53fffffff"),
                (x"fffffffe94eb9cd739ad6b5ad6b5ce777bdefbbd633fffffff"),
                (x"fffffffe94eb9cd739ad6b5ad6b5ce777bdefbbd633fffffff"),
                (x"fffffffe94739ce6b5cd6b5ae777bded3bdef523ef7fffffff"),
                (x"ffffffd3bd739ce739ae739dded3bdf77bdedeecffffffffff"),
                (x"ffffffd3bd739ce739ceef7b4efbdeef6f7bdd20ffffffffff"),
                (x"ffffffd3bdeb9ce73bb4a77bdef7bdbdef7bdd8cffffffffff"),
                (x"ffffff8294a77b4a53bda77bdba58c632f7bdd9fffffffffff"),
                (x"ffffff8294a77b4a53bda77bdba58c632f7bdd9fffffffffff"),
                (x"fffffffc00f5294a53bde8c77ba4a5002f7bdc1fffffffffff"),
                (x"ffffffffffa77bda52891a537ba484002f7bdc1fffffffffff"),
                (x"ffffffffffa33b4a52971a537bdc84ef6f7bdc1fffffffffff"),
                (x"ffffffffffa769def69462537bdc84f7af7bdc1fffffffffff"),
                (x"ffffffffffa769def69462537bdc84f7af7bdc1fffffffffff"),
                (x"fffffffffffd29d633b4a2537bdef7bdef7bdc1fffffffffff"),
                (x"ffffffffffffff4ef694a3189bdef7bdef7ba41fffffffffff"),
                (x"fffffffffffffffa5294a528c4def7bdee9483ffffffffffff"),
                (x"fffffffffffffffef7beef7b46318c6300007fffffffffffff"),
                (x"fffffffffffffffef7beef7b46318c6300007fffffffffffff"),
                (x"ffffffffffffffdef7def529ded000003fffffffffffffffff"),
                (x"ffffffffffffffdf7bdef529df7694a53bffffffffffffffff"),
                (x"ffffffffffffffda50b4077b4f7a94ed3bffffffffffffffff"),
                (x"fffffffffffffe06312c05294ef4006d01ffffffffffffffff"),
                (x"fffffffffffffe06312c05294ef4006d01ffffffffffffffff"),
                (x"fffffffffffffe0bdef767bdebdc006801ffffffffffffffff"),
                (x"fffffffffffffe04a6f74fbdebdc00a001ffffffffffffffff"),
                (x"ffffffffffffffdef5374d294ba7bdef41ffffffffffffffff"),
                (x"ffffffffffffffda53a0a529400294e03bffffffffffffffff"),
                (x"ffffffffffffffda53a0a529400294e03bffffffffffffffff"),
                (x"ffffffffffffffda529df7bdded294e741ffffffffffffffff"),
                (x"fffffffffffffe0a529df7bdda53bde741ffffffffffffffff"),
                (x"fffffffffffffff0001cef7ae73bbde7ffffffffffffffffff"),
                (x"ffffffffffffffffffe00739def000ffffffffffffffffffff"),
                (x"ffffffffffffffffffe00739def000ffffffffffffffffffff"),
                (x"ffffffffffffffffffff00014a0000ffffffffffffffffffff"),

                -- 5_character_0_2
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffe9d739cd6b5ad6b5ad6bbbded29fffffffffff"),
                (x"ffffffffffa75cd6b5ad6b5ad6b5ad739ce777bda53fffffff"),
                (x"ffffffffffa75cd6b5ad6b5ad6b5ad739ce777bda53fffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ce775ce73bbdef69ffffff"),
                (x"ffffffd3bd739ceef7bdf7bdef7bdeed294a77bdef7b4fffff"),
                (x"ffffffd3bd73a94ef7b4ef7bdef7bded294a529def7b4fffff"),
                (x"ffffffd3bd73a94ef7b4ef7bdef7bded294a529def7b4fffff"),
                (x"ffffffd294ef7b4ef7bdeb1831b18cef7bded29def7b4fffff"),
                (x"ffffff8294ed3bd6319d4b18318d8c4f59def7b4ef680fffff"),
                (x"fffffffc00ef7bd4a6f7bdee91a6f7bdeec677bdef41ffffff"),
                (x"fffffffe940307dbdef7bdef7bdef7bdef7bf47d0029ffffff"),
                (x"fffffffe9460d9d632f7bdef7bdef7bdeec67583ef69ffffff"),
                (x"fffffffe9460d9d632f7bdef7bdef7bdeec67583ef69ffffff"),
                (x"ffffffffffeb3a94a6f7bdef7bdef7bdee94a68cef7fffffff"),
                (x"ffffffffffa33a9bdd8c65ef7bdef7631894a68ca53fffffff"),
                (x"ffffffffff053a9bdca005ef7bdef7000b7ba694003fffffff"),
                (x"ffffffffff05e89bdc8005ef7bdef700097ba697003fffffff"),
                (x"ffffffffff05e89bdc8005ef7bdef700097ba697003fffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"ffffffffffffc0cbdc9ef5ef7bdef7f7897bb01fffffffffff"),
                (x"fffffffffffffa04a6f7bdef7bdef7bdee9483bfffffffffff"),
                (x"ffffffffffed3b463137bdef7bdef7bdd2c653b4ef7fffffff"),
                (x"ffffffffffed3b463137bdef7bdef7bdd2c653b4ef7fffffff"),
                (x"ffffffffbdefbbda53ac4a537bdd294b3b4a77beef7bffffff"),
                (x"fffffff7bdf7bb4a53bda318c6318ca77b4a53bef7bbdfffff"),
                (x"ffffff8000a5294a53bef5280a0294f7bb4a5294a5000fffff"),
                (x"fffff626f7bb29da53def77ada37bdf7bd4a768cbdee967fff"),
                (x"fffff626f7bb29da53def77ada37bdf7bd4a768cbdee967fff"),
                (x"fffff6258cf5280a53bef000deb400f7bb4a0294f798967fff"),
                (x"ffffff83dea2580ef69df001405000f769de8189a53c0fffff"),
                (x"ffffff8294bdd2ca5294a77bdef7bda5294a3137bde80fffff"),
                (x"fffffffc00bdd20a53bde8014ed000ef7b4a0137bdc1ffffff"),
                (x"fffffffc00bdd20a53bde8014ed000ef7b4a0137bdc1ffffff"),
                (x"ffffffffff00000a53bef001d77400f7bb4a0000003fffffff"),
                (x"fffffffffffffffef7bdeb9dce71ceef7bdeffffffffffffff"),
                (x"fffffffffffffffe73ad6b9dd075ce6b7bce7fffffffffffff"),
                (x"fffffffffffffff003ae777bd077bd73ba007fffffffffffff"),
                (x"fffffffffffffff003ae777bd077bd73ba007fffffffffffff"),
                (x"fffffffffffffffffe94a5294fd294a529ffffffffffffffff"),

                -- 5_character_0_3
                (x"fffffffffffffbdef7bdef7bda53ffffffffffffffffffffff"),
                (x"ffffffffffa75ce6b5ad6b5ae777bda53fffffffffffffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad777b4a77ffffffffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad777b4a77ffffffffffff"),
                (x"fffffffe94735ad6b5ad6b5ad6b5ad6b5ddef69fffffffffff"),
                (x"fffffffe94a77ae6b5ad6b5ad6b5ad6b5ae73bb4ffffffffff"),
                (x"fffffffd8cef7ddef7ae735ad6b5ad6b5cd6b9dda53fffffff"),
                (x"fffffffd8cef7ddef7ae735ad6b5ad6b5cd6b9dda53fffffff"),
                (x"ffffffffbd1a7bdef69def7ae735ad6b9ae739cea53fffffff"),
                (x"ffffffffff65efdef7beed29deb9ce735ce739ceef69ffffff"),
                (x"ffffffffff026f7bdfbdefbdda77bd739ce739ceef69ffffff"),
                (x"ffffffffff632f7bdef7bf7bdef694a75ce739ddef69ffffff"),
                (x"fffffffffffb2f7bdd8c62537ef694ef694a77b4a501ffffff"),
                (x"fffffffffffb2f7bdd8c62537ef694ef694a77b4a501ffffff"),
                (x"fffffffffff82f7bdc002a537b8c6367694a529e003fffffff"),
                (x"fffffffffff82f7bdc0022537ba4634d29def7b4ffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba463bd294a7594ffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba58ca53bded3b4ffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba58ca53bded3b4ffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694a759ded29fffffffffff"),
                (x"fffffffffff8137bdef7bdef74b294a53b4a7fffffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a529ffffffffffffffff"),
                (x"fffffffffffffe00018c6318ca77bdf77bffffffffffffffff"),
                (x"fffffffffffffe00018c6318ca77bdf77bffffffffffffffff"),
                (x"fffffffffffffffffc000529ded3def7bbdeffffffffffffff"),
                (x"fffffffffffffffef694a77beed3def7bddeffffffffffffff"),
                (x"fffffffffffffffef69da7bdea7400a769deffffffffffffff"),
                (x"fffffffffffffff0028d077bda50006258007fffffffffffff"),
                (x"fffffffffffffff0028d077bda50006258007fffffffffffff"),
                (x"fffffffffffffff0000d05ef7f798cbdee007fffffffffffff"),
                (x"fffffffffffffff0001405ef7f7929bdd2007fffffffffffff"),
                (x"fffffffffffffff003bdea537a5129ba7bdeffffffffffffff"),
                (x"fffffffffffffffef41ca0000a52940769deffffffffffffff"),
                (x"fffffffffffffffef41ca0000a52940769deffffffffffffff"),
                (x"fffffffffffffff003bca529defbdeed29deffffffffffffff"),
                (x"fffffffffffffff003bced294efbdeed28007fffffffffffff"),
                (x"fffffffffffffffffffceb9ce777bde001ffffffffffffffff"),
                (x"ffffffffffffffffffff0739def00007ffffffffffffffffff"),
                (x"ffffffffffffffffffff0739def00007ffffffffffffffffff"),
                (x"ffffffffffffffffffff00014a0000ffffffffffffffffffff"),

                -- 5_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffe9def5ce739ce739ce739ddef69fffffffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b9ae739dda53fffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad6b5cd6b9ceef69ffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad6b5cd6b9ceef69ffffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae739ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ae735ce739d4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4fffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae735cd73bb4fffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae735cd73bb4fffff"),
                (x"ffffffd3bdeb9cd6b5ad6b5ad6b5ad6b5ad6b9aeef7b4fffff"),
                (x"ffffffd294ef7ae739cd6b5ad6b5ad6b5ae73bbdef694fffff"),
                (x"fffffffe94ef7bdef7ae739ce739ce73bbdef7bdef69ffffff"),
                (x"ffffffffffa53bdef7bdef7bdef7bdef7bdef7bda53bffffff"),
                (x"ffffffffffa53bdef7bdef7bdef7bdef7bdef7bda53bffffff"),
                (x"ffffffffffef694a53bdef7bdef7bdef7b4a529def7fffffff"),
                (x"ffffffffffff7b4a5294a77bdef7bda5294a53a0ffffffffff"),
                (x"ffffffffffffc1def7b4ef7bdef7bded3bdef41fffffffffff"),
                (x"fffffffffffffe0a53aca3194ef7bdef594a03ffffffffffff"),
                (x"fffffffffffffe0a53aca3194ef7bdef594a03ffffffffffff"),
                (x"fffffffffffd29da529da77b4ed3bda5294a529fffffffffff"),
                (x"ffffffffffa53deef694a5294a5294053bef7a94ffffffffff"),
                (x"ffffffffff07bdea53beed294a5000a53bef7bd4ffffffffff"),
                (x"ffffffffff483dda53bef4e619fbdeef7bef5000a53fffffff"),
                (x"ffffffffff483dda53bef4e619fbdeef7bef5000a53fffffff"),
                (x"ffffffffff65c00a53bef7bdef7bdef53a005eeca53fffffff"),
                (x"ffffffffff03180a529df04330fbdeed017bdee9633fffffff"),
                (x"fffffffffff8014a5294a77bded294a50094dee9633fffffff"),
                (x"ffffffffffffff4a529defbdeefbdeef68c62520ffffffffff"),
                (x"ffffffffffffff4a529defbdeefbdeef68c62520ffffffffff"),
                (x"ffffffffffffff4a529df7bdeef7deed294a001fffffffffff"),
                (x"fffffffffffffffe739ceb9ceef39ce700007fffffffffffff"),
                (x"fffffffffffffffffc1d735ae7779ce03fffffffffffffffff"),
                (x"fffffffffffffffffffc777bde839ce7ffffffffffffffffff"),
                (x"fffffffffffffffffffc777bde839ce7ffffffffffffffffff"),
                (x"ffffffffffffffffffff00000003ffffffffffffffffffffff"),

                -- 5_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffd294ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffffffd294ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffe94ef7ae735ad6b5ae73bb4ffffffffff"),
                (x"ffffffffffffff4ef7ae6b5ad6b5ad6b5ad6b5dda53fffffff"),
                (x"fffffffffffd3bd739ad6b5ad6b5ad6b5ad6b5aea53fffffff"),
                (x"fffffffffffd3bd739ad6b5ad6b5ad6b5ad6b5aea53fffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b5ae777b4a53fffffff"),
                (x"fffffffe94eb9cd739ad6b5ad6b5ce777bdefbbd633fffffff"),
                (x"fffffffe94739ce6b5cd6b5ae777bded3bdef523ef7fffffff"),
                (x"ffffffd3bd739ce739ae739dded3bdf77bdedeecffffffffff"),
                (x"ffffffd3bd739ce739ceef7b4efbbdef6f7bdd20ffffffffff"),
                (x"ffffffd3bd739ce739ceef7b4efbbdef6f7bdd20ffffffffff"),
                (x"ffffffd3bdeb9ce73bb4a77bdef6f7bdef7bdd8cffffffffff"),
                (x"ffffff8294a77b4a53bda77bdba58c632f7bdd9fffffffffff"),
                (x"fffffffc00f5294a53bd18c77ba4a5002f7bdc1fffffffffff"),
                (x"ffffffffff077bda52891a537ba484002f7bdc1fffffffffff"),
                (x"ffffffffff077bda52891a537ba484002f7bdc1fffffffffff"),
                (x"ffffffffffa33b4a52971a537bdc84ef6f7bdc1fffffffffff"),
                (x"ffffffffffa769def69462537bdc84f7af7bdc1fffffffffff"),
                (x"fffffffffffd29d633b4a2537bdef7bdef7bdc1fffffffffff"),
                (x"ffffffffffffff4ef694a3189bdef7bdef7ba41fffffffffff"),
                (x"ffffffffffffff4ef694a3189bdef7bdef7ba41fffffffffff"),
                (x"fffffffffffffffa5294a528c4def7bdee9483ffffffffffff"),
                (x"ffffffffffffffffffbded29d6318c6300007fffffffffffff"),
                (x"fffffffffffffffef7bef77b4a0000003fffffffffffffffff"),
                (x"fffffffffffffff003def7bdda7400e83bffffffffffffffff"),
                (x"fffffffffffffff003def7bdda7400e83bffffffffffffffff"),
                (x"fffffffffffffff003bda77a0ef400a03bffffffffffffffff"),
                (x"fffffffffffffe0ef41463194a26f7483bffffffffffffffff"),
                (x"fffffffffffffe0a500cbdef4f26f7b801ffffffffffffffff"),
                (x"ffffffffffffffda5289bdee9f5129b83bffffffffffffffff"),
                (x"ffffffffffffffda5289bdee9f5129b83bffffffffffffffff"),
                (x"ffffffffffffc14ef6804def7f7a94077bffffffffffffffff"),
                (x"ffffffffffffc14a53bd00000a039ca53bffffffffffffffff"),
                (x"fffffffffffffe0ef694a77bd073bdef7fffffffffffffffff"),
                (x"fffffffffffffe0e73bd739dd073bde801ffffffffffffffff"),
                (x"fffffffffffffe0e73bd739dd073bde801ffffffffffffffff"),
                (x"fffffffffffffff0000000000003ffffffffffffffffffffff"),

                -- 5_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffe9d739cd6b5ad6b5ad6bbbded29fffffffffff"),
                (x"ffffffffffffe9d739cd6b5ad6b5ad6bbbded29fffffffffff"),
                (x"ffffffffffa75cd6b5ad6b5ad6b5ad739ce777bda53fffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ce775ce73bbdef69ffffff"),
                (x"ffffffd3bd739ceef7bdf7bdef7bdeed294a77bdef7b4fffff"),
                (x"ffffffd3bd739ceef7bdf7bdef7bdeed294a77bdef7b4fffff"),
                (x"ffffffd3bd73a94ef7b4ef7bdef7bded294a529def7b4fffff"),
                (x"ffffffd294ef7b4ef7bdeb1831b18cef7bded29def7b4fffff"),
                (x"ffffff8294ed3bd6319d4b18318d8c4f59def7b4ef680fffff"),
                (x"fffffffc00ef7bd4a6f7bdee91a6f7bdeec677bdef41ffffff"),
                (x"fffffffe940307dbdef7bdef7bdef7bdef7bf47d0029ffffff"),
                (x"fffffffe940307dbdef7bdef7bdef7bdef7bf47d0029ffffff"),
                (x"fffffffe9460d9d632f7bdef7bdef7bdeec67583ef69ffffff"),
                (x"ffffffffffeb3a94a6f7bdef7bdef7bdee94a68cef7fffffff"),
                (x"ffffffffffa33a9bdd8c65ef7bdef7631894a68ca53fffffff"),
                (x"ffffffffff053a9bdca005ef7bdef7000b7ba694003fffffff"),
                (x"ffffffffff053a9bdca005ef7bdef7000b7ba694003fffffff"),
                (x"ffffffffff05e89bdc8005ef7bdef700097ba697003fffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"ffffffffffffc0cbdc9ef5ef7bdef7f7897bb01fffffffffff"),
                (x"fffffffffffffa04a6f7bdef7bdef7bdee9483ffffffffffff"),
                (x"fffffffffffffa04a6f7bdef7bdef7bdee9483ffffffffffff"),
                (x"ffffffffffff69d63137bdef7bdef7bdd2c6769def7fffffff"),
                (x"ffffffffffed3dda528c4a537bdd294b3b4a77dda53bffffff"),
                (x"fffffffc00a77bda53bda1ce739ce7a7694a7bdeef7bffffff"),
                (x"fffffffd8c653b4a53bef5280a0294f7a9de829d0029dfffff"),
                (x"fffffffd8c653b4a53bef5280a0294f7a9de829d0029dfffff"),
                (x"fffffff9294b014a53def77adeb7bdf7a80001974a41dfffff"),
                (x"ffffffd3def781da53def528deb694f780c652944a59ffffff"),
                (x"ffffffb294a5000ef69df001405000ef597ba694003fffffff"),
                (x"ffffffb129bb01da53b4a529def7bdef597bdd34003fffffff"),
                (x"ffffffb129bb01da53b4a529def7bdef597bdd34003fffffff"),
                (x"ffffff8129483fda53def001d77400a50094dd20ffffffffff"),
                (x"fffffffc00003e0ef694a001de7400ef7800001fffffffffff"),
                (x"fffffffffffffff003bd735aee83bdef3fffffffffffffffff"),
                (x"ffffffffffffffffff9d735aee83bde83fffffffffffffffff"),
                (x"ffffffffffffffffff9d735aee83bde83fffffffffffffffff"),
                (x"ffffffffffffffffffe00000000000ffffffffffffffffffff"),

                -- 5_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffbdef7bdef7bda53ffffffffffffffffffffff"),
                (x"fffffffffffffbdef7bdef7bda53ffffffffffffffffffffff"),
                (x"ffffffffffa75ce6b5ad6b5ae777bda53fffffffffffffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad777b4a77ffffffffffff"),
                (x"fffffffe94735ad6b5ad6b5ad6b5ad6b5ddef69fffffffffff"),
                (x"fffffffe94735ad6b5ad6b5ad6b5ad6b5ddef69fffffffffff"),
                (x"fffffffe94a77ad6b5ad6b5ad6b5ad6b5ae73bb4ffffffffff"),
                (x"fffffffd8cef7ddef7ae735ad6b5ad6b5cd6b9dda53fffffff"),
                (x"ffffffffbd1a7bdef69def7ae735ad6b9ae739cea53fffffff"),
                (x"ffffffffff65efdef7beed29deb9ce735ce739ceef69ffffff"),
                (x"ffffffffff026f7bdefdefbdda77bd739ce739ceef69ffffff"),
                (x"ffffffffff026f7bdefdefbdda77bd739ce739ceef69ffffff"),
                (x"ffffffffff632f7bdef7bf7bdef694a75ce739ddef69ffffff"),
                (x"fffffffffffb2f7bdd8c62537ef694ef694a77b4a501ffffff"),
                (x"fffffffffff82f7bdc002a537b8c63ef694a529e003fffffff"),
                (x"fffffffffff82f7bdc0022537ba4634d3bdef7a0ffffffffff"),
                (x"fffffffffff82f7bdc0022537ba4634d3bdef7a0ffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba463bd294a7594ffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba58ca53bded3b4ffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694a759ded29fffffffffff"),
                (x"fffffffffff8137bdef7bdef74b294a53b4a7fffffffffffff"),
                (x"fffffffffff8137bdef7bdef74b294a53b4a7fffffffffffff"),
                (x"ffffffffffffc09bdef7bdee965294a529ffffffffffffffff"),
                (x"fffffffffffffe00018c6318ced3bdef7fffffffffffffffff"),
                (x"fffffffffffffffffc0000014a77def77bffffffffffffffff"),
                (x"fffffffffffffffef41d077b4efbdef781ffffffffffffffff"),
                (x"fffffffffffffffef41d077b4efbdef781ffffffffffffffff"),
                (x"fffffffffffffffef414077bd07694ef41ffffffffffffffff"),
                (x"fffffffffffffffef409ba534a318ca03a007fffffffffffff"),
                (x"fffffffffffffff00017ba53ea5ef76028007fffffffffffff"),
                (x"fffffffffffffffef4174d29e4def74d29deffffffffffffff"),
                (x"fffffffffffffffef4174d29e4def74d29deffffffffffffff"),
                (x"fffffffffffffffef7a0a7bdebdd29053b4a03ffffffffffff"),
                (x"fffffffffffffffef694e001400000ef694a03ffffffffffff"),
                (x"fffffffffffffffffc1def380ef694a53a007fffffffffffff"),
                (x"fffffffffffffff0001def380eb9ceef78007fffffffffffff"),
                (x"fffffffffffffff0001def380eb9ceef78007fffffffffffff"),
                (x"fffffffffffffffffffffffe0000000001ffffffffffffffff"),

                -- 5_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffe9def5ce739ce739ce739ddef69fffffffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b9ae739dda53fffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad6b5cd6b9ceef69ffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad6b5cd6b9ceef69ffffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae739ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce73bb4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ae735ce739d4fffff"),
                (x"ffffffd1ce6b5ad6b5ad6b5ad6b5ad6b5ad6b9ce739d4fffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae735cd73bb4fffff"),
                (x"ffffffd3bd735ad6b5ad6b5ad6b5ad6b5ae735cd73bb4fffff"),
                (x"ffffffd3bdeb9cd6b5ad6b5ad6b5ad6b5ad6b9aeef7b4fffff"),
                (x"ffffffd294ef7ae739cd6b5ad6b5ad6b5ae73bbdef694fffff"),
                (x"fffffffe94ef7bdef7ae739ce739ce73bbdef7bdef69ffffff"),
                (x"ffffffffffa53bdef7bdef7bdef7bdef7bdef7bda53bffffff"),
                (x"ffffffffffa53bdef7bdef7bdef7bdef7bdef7bda53bffffff"),
                (x"ffffffffffef694a53bdef7bdef7bdef7b4a529def7fffffff"),
                (x"ffffffffffff7b4a5294a77bdef7bda5294a53bdffffffffff"),
                (x"ffffffffffffc14ef7b4ef7bdef7bded3bdef41fffffffffff"),
                (x"fffffffffffffe0a53aca77bdef7bdef594a03ffffffffffff"),
                (x"fffffffffffffe0a53aca77bdef7bdef594a03ffffffffffff"),
                (x"ffffffffffffe94a529da77b4ed3bda5294a7694ffffffffff"),
                (x"fffffffffffd29ef7bb405294a5294a529defbd4a53fffffff"),
                (x"fffffffffffd3def7bb4a0014a5294efbb4a7bde003fffffff"),
                (x"ffffffffffa0014f7bbdefbde98673f7bb4a77c04a7fffffff"),
                (x"ffffffffffa0014f7bbdefbde98673f7bb4a77c04a7fffffff"),
                (x"ffffffffffa32f7003b4f7bdef7bdef7bb4a0017633fffffff"),
                (x"ffffffffff626f7bdc14efbde0cc21f7694a018c003fffffff"),
                (x"ffffffffff626f74a414a5294ef7bda5294a5000ffffffffff"),
                (x"fffffffffff81296329defbdeefbdeef694a53ffffffffffff"),
                (x"fffffffffff81296329defbdeefbdeef694a53ffffffffffff"),
                (x"ffffffffffffc00a5294efbddefbdef7694a53ffffffffffff"),
                (x"fffffffffffffff0001ce739ceb9ceef39ce7fffffffffffff"),
                (x"ffffffffffffffffffe0e739d739ad7741ffffffffffffffff"),
                (x"ffffffffffffffffffffe7380ef7bd773fffffffffffffffff"),
                (x"ffffffffffffffffffffe7380ef7bd773fffffffffffffffff"),
                (x"fffffffffffffffffffffffe000000e7ffffffffffffffffff"),

                -- 5_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffd294ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffffffd294ef7bdef7bdef7ffffffffffff"),
                (x"fffffffffffffffffe94ef7ae735ad6b5ae73bb4ffffffffff"),
                (x"ffffffffffffff4ef7ae6b5ad6b5ad6b5ad6b5dda53fffffff"),
                (x"fffffffffffd3bd739ad6b5ad6b5ad6b5ad6b5aea53fffffff"),
                (x"fffffffffffd3bd739ad6b5ad6b5ad6b5ad6b5aea53fffffff"),
                (x"ffffffffffa75ce6b5ad6b5ad6b5ad6b5ae777b4a53fffffff"),
                (x"fffffffe94eb9cd739ad6b5ad6b5ce777bdefbbd633fffffff"),
                (x"fffffffe94739ce6b5cd6b5ae777bded3bdef5237bffffffff"),
                (x"ffffffd3bd739ce739ae739dded3bdf77bdedeecffffffffff"),
                (x"ffffffd3bd739ce739ceef7b4efbdeef6f7bdd20ffffffffff"),
                (x"ffffffd3bd739ce739ceef7b4efbdeef6f7bdd20ffffffffff"),
                (x"ffffffd3bdeb9ce73bb4a77bdef7bdbdef7bdd8cffffffffff"),
                (x"ffffff8294a77b4a53bda77bdba58c632f7bdd9fffffffffff"),
                (x"fffffffc00f5294a53bde8c77ba4a5002f7bdc1fffffffffff"),
                (x"ffffffffff077bdef6891a537ba484002f7bdc1fffffffffff"),
                (x"ffffffffff077bdef6891a537ba484002f7bdc1fffffffffff"),
                (x"ffffffffffa33b4a52971a537bdc84ef6f7bdc1fffffffffff"),
                (x"ffffffffffa769def69462537bdc84f7af7bdc1fffffffffff"),
                (x"fffffffffffd29d633b4a2537bdef7bdef7bdc1fffffffffff"),
                (x"ffffffffffffff4ef694a3189bdef7bdef7ba41fffffffffff"),
                (x"ffffffffffffff4ef694a3189bdef7bdef7ba41fffffffffff"),
                (x"fffffffffffffffa5294ed28c4def7bdee9483ffffffffffff"),
                (x"ffffffffffffffdef7dda77b439ce739c0007fffffffffffff"),
                (x"fffffffffffffbdf7bdeefbdee83bd0741ffffffffffffffff"),
                (x"ffffffffffffe94ef7bea7bdef03bd07414a7fffffffffffff"),
                (x"ffffffffffffe94ef7bea7bdef03bd07414a7fffffffffffff"),
                (x"ffffffffffffc0063194ef7bef51ada340c67fffffffffffff"),
                (x"ffffffffffffc094a520ed29df51ada76894b3ffffffffffff"),
                (x"ffffffffffffc09bdd3ef529ded3bda5009483ffffffffffff"),
                (x"ffffffffffffc0c4a69ea2529a5294ef40007fffffffffffff"),
                (x"ffffffffffffc0c4a69ea2529a5294ef40007fffffffffffff"),
                (x"fffffffffffffe06329ea5ef7077dea77bffffffffffffffff"),
                (x"ffffffffffffffdef414a5ef7077bda77bffffffffffffffff"),
                (x"fffffffffffffe0003bda5294a5294ef01ffffffffffffffff"),
                (x"fffffffffffffffe739ce739deb800073fffffffffffffffff"),
                (x"fffffffffffffffe739ce739deb800073fffffffffffffffff"),
                (x"fffffffffffffff0039cf80000039ce001ffffffffffffffff"),

                -- 5_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffa5294ef7bdef7bded294a7fffffffffffff"),
                (x"ffffffffffffe9d739cd6b5ad6b5ad6bbbded29fffffffffff"),
                (x"ffffffffffffe9d739cd6b5ad6b5ad6bbbded29fffffffffff"),
                (x"ffffffffffa75cd6b5ad6b5ad6b5ad739ce777bda53fffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ce775ce73bbdef69ffffff"),
                (x"ffffffd3bd739ceef7bdf7bdef7bdeed294a77bdef7b4fffff"),
                (x"ffffffd3bd739ceef7bdf7bdef7bdeed294a77bdef7b4fffff"),
                (x"ffffffd3bd73a94ef7b4ef7bdef7bded294a529def7b4fffff"),
                (x"ffffffd294ef7b4ef7bdeb1831b18cef7bded29def7b4fffff"),
                (x"ffffff8294ed3bd6319d4b18318d8c4f59def7b4ef680fffff"),
                (x"fffffffc00ef7bd4a6f7bdee91a6f7bdeec677bdef41ffffff"),
                (x"fffffffe940307dbdef7bdef7bdef7bdef7bf47d0029ffffff"),
                (x"fffffffe940307dbdef7bdef7bdef7bdef7bf47d0029ffffff"),
                (x"fffffffe9460d9d632f7bdef7bdef7bdeec67583ef69ffffff"),
                (x"ffffffffffeb3a94a6f7bdef7bdef7bdee94a68cef7fffffff"),
                (x"ffffffffffa33a9bdd8c65ef7bdef7631894a68ca53fffffff"),
                (x"ffffffffff053a9bdca005ef7bdef7000b7ba694003fffffff"),
                (x"ffffffffff053a9bdca005ef7bdef7000b7ba694003fffffff"),
                (x"ffffffffff05e89bdc8005ef7bdef700097ba697003fffffff"),
                (x"fffffffffff8009bdc9dedef7bdef7ef497ba400ffffffffff"),
                (x"ffffffffffffc0cbdc9ef5ef7bdef7f7897bb01fffffffffff"),
                (x"fffffffffffffe04a6f7bdef7bdef7bdee9483bfffffffffff"),
                (x"fffffffffffffe04a6f7bdef7bdef7bdee9483bfffffffffff"),
                (x"ffffffffffef69d63137bdef7bdef7bdd2c6769dffffffffff"),
                (x"ffffffffbda77dda53ac4a537bdd294b294a77d4ef7fffffff"),
                (x"ffffffffbdefbdea529da1ce739ce7a77b4a77bda501ffffff"),
                (x"fffffff69407680ef69ef5280a0294f7bb4a53b46319ffffff"),
                (x"fffffff69407680ef69ef5280a0294f7bb4a53b46319ffffff"),
                (x"fffffff4004dd800029ef77adeb7bdf7bd4a500c4a52cfffff"),
                (x"fffffffd8c4d2946301ef528deb694f7bd4a741ef7bccfffff"),
                (x"ffffffffff05289bdd9de801405000f769de8014a529ffffff"),
                (x"ffffffffff05137bdd9def7bdef694a53b4a740cbdd3ffffff"),
                (x"ffffffffff05137bdd9def7bdef694a53b4a740cbdd3ffffff"),
                (x"fffffffffff81374a414a001d77400f7bd4a77e04a53ffffff"),
                (x"ffffffffffffc000039de801de7400a529de83e00001ffffff"),
                (x"fffffffffffffffffffcef7a0eb9ad777a007fffffffffffff"),
                (x"ffffffffffffffffffe0ef7a0eb9ad7779ffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7a0eb9ad7779ffffffffffffffff"),
                (x"fffffffffffffffffffff8000e0000003fffffffffffffffff"),

                -- 5_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffbdef7bdef7bda53ffffffffffffffffffffff"),
                (x"fffffffffffffbdef7bdef7bda53ffffffffffffffffffffff"),
                (x"ffffffffffa75ce6b5ad6b5ae777bda53fffffffffffffffff"),
                (x"fffffffe94eb9ad6b5ad6b5ad6b5ad777b4a7fffffffffffff"),
                (x"fffffffe94735ad6b5ad6b5ad6b5ad6b5ddef69fffffffffff"),
                (x"fffffffe94735ad6b5ad6b5ad6b5ad6b5ddef69fffffffffff"),
                (x"fffffffe94a77ae6b5ad6b5ad6b5ad6b5ae73bb4ffffffffff"),
                (x"fffffffd8cef7ddef7ae735ad6b5ad6b5cd6b9dda53fffffff"),
                (x"ffffffffbd1a7bdef69def7ae735ad6b9ae739cea53fffffff"),
                (x"ffffffffff65efdef7beed29deb9ce735ce739ceef69ffffff"),
                (x"ffffffffff026f7bdfbdefbdda77bd739ce739ceef69ffffff"),
                (x"ffffffffff026f7bdfbdefbdda77bd739ce739ceef69ffffff"),
                (x"ffffffffff632f7bdef7bf7bdef694a75ce739ddef69ffffff"),
                (x"fffffffffffb2f7bdd8c62537ef694ef694a77b4a501ffffff"),
                (x"fffffffffff82f7bdc002a537b8c63ef694a529e003fffffff"),
                (x"fffffffffff82f7bdc0022537ba4634d29def7a0ffffffffff"),
                (x"fffffffffff82f7bdc0022537ba4634d29def7a0ffffffffff"),
                (x"fffffffffff82f7bdfbd25ef7ba463bd294a7594ffffffffff"),
                (x"fffffffffff82f7bdfde25ef7ba58ca53bded3b4ffffffffff"),
                (x"fffffffffff82f7bdef7bdef7ba694a759ded29fffffffffff"),
                (x"fffffffffff8137bdef7bdef74b294a53b4a7fffffffffffff"),
                (x"fffffffffff8137bdef7bdef74b294a53b4a7fffffffffffff"),
                (x"ffffffffffffc09bdef7bdee9653bda529ffffffffffffffff"),
                (x"fffffffffffffe00018c6318ca7694efbbdeffffffffffffff"),
                (x"fffffffffffffff003a0e801df7bbdf7bddef7ffffffffffff"),
                (x"ffffffffffffff4003a0e801ef7a94f77b4a53ffffffffffff"),
                (x"ffffffffffffff4003a0e801ef7a94f77b4a53ffffffffffff"),
                (x"fffffffffffffec001b46d29ef77bda3180003ffffffffffff"),
                (x"ffffffffffffd89a53b46d29eed3bd02529483ffffffffffff"),
                (x"ffffffffffffc0900294ed29ded3def26e9483ffffffffffff"),
                (x"fffffffffffffe0003bda52944a694f512c603ffffffffffff"),
                (x"fffffffffffffe0003bda52944a694f512c603ffffffffffff"),
                (x"fffffffffffffffef7b4f77a0bde94f518007fffffffffffff"),
                (x"fffffffffffffffef7b4ef7a0bde94a03bdeffffffffffffff"),
                (x"fffffffffffffff0039da5294a5294ef40007fffffffffffff"),
                (x"ffffffffffffffffff8e739ddef39ce739ffffffffffffffff"),
                (x"ffffffffffffffffff8e739ddef39ce739ffffffffffffffff"),
                (x"fffffffffffffff0000000000003ffe701ffffffffffffffff"),

                -- 6_character_0_0
                (x"fffffffffffffffffd8cef7bdef7bded29ffffffffffffffff"),
                (x"ffffffffffffff4a53bef0c7eefbdef77ac633ffffffffffff"),
                (x"fffffffffffd3bef7bddf0c63f0fdef769def7b4ffffffffff"),
                (x"fffffffffffd3bef7bddf0c63f0fdef769def7b4ffffffffff"),
                (x"ffffffffffa77c318fdef0c6318fdef53b4a77dda53fffffff"),
                (x"ffffffffffa53be18c7eefbc318fdeed29defbb4a53fffffff"),
                (x"fffffffc00ef69df787eefbc3f0fdeed3bef769def69ffffff"),
                (x"fffffffc00ef69df787eefbc3f0fdeed3bef769def69ffffff"),
                (x"fffffffc00a7bb4ef7bef77bee8fbda53bded3bea501ffffff"),
                (x"fffffffc00a77dda529df77beefbbda77b4a03dda501ffffff"),
                (x"fffffffc00ed3beef694ef7bda7694a7680053b4a501ffffff"),
                (x"fffffffc00a7694ef694a529da7694a5294a50140001ffffff"),
                (x"ffffffffff077bda5294a5294a5294a5294a0294003fffffff"),
                (x"ffffffffff077bda5294a5294a5294a5294a0294003fffffff"),
                (x"ffffffffff053bdef694ed294a5294a528005280003fffffff"),
                (x"ffffffffff053bdef7b4ed294a5294a5294a5000003fffffff"),
                (x"ffffffffff053beef7bdef7b4a7694a5294a0280003fffffff"),
                (x"ffffffffffa77bea53bdf77b4ef694a7694a5294003fffffff"),
                (x"ffffffffffa77bea53bdf77b4ef694a7694a5294003fffffff"),
                (x"ffffffffffa77bea53bdf77bdefbbda7694a5014003fffffff"),
                (x"ffffffffffefbbdf7a9df77b4efbbda53b4a5014003fffffff"),
                (x"ffffffffffefa9df781df7bd4f7bbda53b4a5014003fffffff"),
                (x"ffffffffffa741df781df7bd4f7bbd053b4a5014003fffffff"),
                (x"ffffffffffa741df781df7bd4f7bbd053b4a5014003fffffff"),
                (x"ffffffffff05014ef414efbc0efa94053a0050004a7fffffff"),
                (x"fffffffcc605000a5014ef7a0a769405280050094a4dffffff"),
                (x"ffffffffde4812000200a5280a500005000001294a7dffffff"),
                (x"fffffffd8c4b19e001e500005000a5281e00798c4a59ffffff"),
                (x"fffffffd8c4b19e001e500005000a5281e00798c4a59ffffff"),
                (x"fffffffc004dd20ef7cf842052961083fdde81374a41ffffff"),
                (x"ffffffffff0000cef7bdf18c6318c6f77bdeb000003fffffff"),
                (x"fffffffffffffe0ef4e77bde7e9def79cfde83ffffffffffff"),
                (x"fffffffffffffffef4e77bde7e9def79cfdeffffffffffffff"),
                (x"fffffffffffffffef4e77bde7e9def79cfdeffffffffffffff"),
                (x"fffffffffffffffef7a739cfdef4e739fbdeffffffffffffff"),
                (x"fffffffffffffff003bdef7bd077bdef7a007fffffffffffff"),
                (x"fffffffffffffff003bd3f7bd077bd3f7a007fffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc0739ce0f80e739c1ffffffffffffffff"),
                (x"fffffffffffffffffc1df77a0f83bdf741ffffffffffffffff"),

                -- 6_character_0_1
                (x"fffffffffffffffffe94ef7bded294ef58c633ffffffffffff"),
                (x"ffffffffffffff4ef7bdefbdef7bdea0fddef694ffffffffff"),
                (x"ffffffffffffe9def694ef7bde8c63f747ef0fbda53fffffff"),
                (x"ffffffffffffe9def694ef7bde8c63f747ef0fbda53fffffff"),
                (x"fffffffffffd3b4ef7bef7bdeef7de1fbc318fbeef7fffffff"),
                (x"ffffffffff0529def7dda5294a53bdf0fc31fba3ef7fffffff"),
                (x"ffffffffff053bdef694a5289bdd29ed3bef769ea53fffffff"),
                (x"ffffffffff053bdef694a5289bdd29ed3bef769ea53fffffff"),
                (x"fffffffc00a5294a53bdea537bdef7bde9def53dffffffffff"),
                (x"fffffffc00a53bdef7b4a2537bdef7bdef7bdeecffffffffff"),
                (x"fffffffc00a529400294a2537bb3bd4def7bdd20ffffffffff"),
                (x"fffffffc00a0000a529dea5374a694ef537bdd94ffffffffff"),
                (x"fffffffc00a7694a53bda77b7ba58ca53b7bde9fffffffffff"),
                (x"fffffffc00a7694a53bda77b7ba58ca53b7bde9fffffffffff"),
                (x"fffffffc00a769da53b4ed297bdca500137bdc1fffffffffff"),
                (x"fffffffc00a769da5294f5297bdc84002f7bdc1fffffffffff"),
                (x"fffffffe94ed3b4a501df5297bdc84e72f7bdc1fffffffffff"),
                (x"fffffffe94e83a0a501df5297bdc8473af7bdc1fffffffffff"),
                (x"fffffffe94e83a0a501df5297bdc8473af7bdc1fffffffffff"),
                (x"fffffffe94a03a0a501df5297bdef7bdef7bdc1fffffffffff"),
                (x"fffffffe94a028000014f5289bdef7bdef7ba41fffffffffff"),
                (x"fffffffc00a000000294eb18c4def7bdee9483ffffffffffff"),
                (x"fffffffc00a0000003c0a319e6318c6300007fffffffffffff"),
                (x"fffffffc00a0000003c0a319e6318c6300007fffffffffffff"),
                (x"fffffffc00a0000f792904206798c6603dffffffffffffffff"),
                (x"fffffffc000001e4a6e9318cff14a5879fef7fffffffffffff"),
                (x"ffffffffff0001ebdee94a526f78a5843def7fffffffffffff"),
                (x"ffffffffffffffebdefef318c003de8421ef7fffffffffffff"),
                (x"ffffffffffffffebdefef318c003de8421ef7fffffffffffff"),
                (x"fffffffffffffe0bdef7ba537ba4002961ef7fffffffffffff"),
                (x"fffffffffffffe0632f7bdef7bdc00815fef7fffffffffffff"),
                (x"fffffffffffffff00137ba537ba40031bdffffffffffffffff"),
                (x"fffffffffffffffffc006318c018c631bfffffffffffffffff"),
                (x"fffffffffffffffffc006318c018c631bfffffffffffffffff"),
                (x"fffffffffffffffffc1def7bde9ce7ed3fffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7bd3bce7a7ffffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7a779fbdffffffffffffffffffff"),
                (x"ffffffffffffffffffff077af7bc00ffffffffffffffffffff"),
                (x"ffffffffffffffffffff077af7bc00ffffffffffffffffffff"),
                (x"ffffffffffffffffffff077be2f800ffffffffffffffffffff"),

                -- 6_character_0_2
                (x"fffffffffffffffffe94ef7bdef7bded29ffffffffffffffff"),
                (x"ffffffffffffff4a53bdf0c7eefbdef77b4a53ffffffffffff"),
                (x"fffffffffffd3beef69ee8c63f0fdeef69def7b4ffffffffff"),
                (x"fffffffffffd3beef69ee8c63f0fdeef69def7b4ffffffffff"),
                (x"ffffffffffa77c3f7bb4f77a318fdeed3b4a77dda53fffffff"),
                (x"ffffffffffa53be18fddf77be1fbbda529defbb4a53fffffff"),
                (x"fffffffc00ef69d18fb4a77bdf77bda53bef769def41ffffff"),
                (x"fffffffc00ef69d18fb4a77bdf77bda53bef769def41ffffff"),
                (x"fffffffc00a7bb4ef5374d29def6944dd34a53bea501ffffff"),
                (x"fffffffc00a77d4bdef7bdee9ea6f7bdef7bd3dda501ffffff"),
                (x"fffffffc00a03b4bdef7bdef7bdef7bdef7bd3b4a501ffffff"),
                (x"fffffffc00a7414633a9bdef7bdef7ba7ac6529da501ffffff"),
                (x"ffffffffffa76894a69dea537bdd29ef6894a41da53fffffff"),
                (x"ffffffffffa76894a69dea537bdd29ef6894a41da53fffffff"),
                (x"ffffffffff077dd4a594a77b7bdfbda51894d3b4003fffffff"),
                (x"ffffffffff077d4bdca002537bdd29000b7bd3d4003fffffff"),
                (x"ffffffffff053d4bdc8005ef7bdef700097bd3d4003fffffff"),
                (x"ffffffffffa53a0bdc9ce5ef7bdef7e7097bd3d4a53fffffff"),
                (x"ffffffffffa53a0bdc9ce5ef7bdef7e7097bd3d4a53fffffff"),
                (x"ffffffffffa03a0bdc8e75ef7bdef773897b83a0a53fffffff"),
                (x"ffffffffffe83a04a6f7bdef7bdef7bdee9483a0ef7fffffff"),
                (x"ffffffffff3028063137bdef7bdef7bdd2c6028031bfffffff"),
                (x"fffffffcc64a6807bccc4a537bdd294b0cf782894a4dffffff"),
                (x"fffffffcc64a6807bccc4a537bdd294b0cf782894a4dffffff"),
                (x"ffffff99294a4c07bde53318c6318c315ef780c94a526fffff"),
                (x"fffff327def25267bde5294be4f8a52c1ef79929f7bc937fff"),
                (x"fffff331294b13e00205294aff3ca5296000792c4a52c37fff"),
                (x"fffff626f7ba58000205294a5294a52960000189bdee967fff"),
                (x"fffff626f7ba58000205294a5294a52960000189bdee967fff"),
                (x"fffff626f74deec000c5294a5294a5294c0032f74a6e967fff"),
                (x"ffffff81294deecef7c6842108421081bddeb2f74a520fffff"),
                (x"fffffffc004dee0ef4fef7bc631bdef78fde82f74a41ffffff"),
                (x"ffffffffff0001fef4e77bdef7bdef79cfdefc00003fffffff"),
                (x"ffffffffff0001fef4e77bdef7bdef79cfdefc00003fffffff"),
                (x"fffffffffffffffa53a779cfda74e779fb4a7fffffffffffff"),
                (x"fffffffffffffff003a739cfd074e739fa007fffffffffffff"),
                (x"fffffffffffffff003af79cfd074e77bfa007fffffffffffff"),
                (x"fffffffffffffffffc1def7a0f83bdef41ffffffffffffffff"),
                (x"fffffffffffffffffc1def7a0f83bdef41ffffffffffffffff"),
                (x"ffffffffffffffffffbdf77a0f83bdf77bffffffffffffffff"),

                -- 6_character_0_3
                (x"ffffffffffffe94a53bda529def7bda53fffffffffffffffff"),
                (x"ffffffffffa53bdf7874f7bdef7bbdef7b4a7fffffffffffff"),
                (x"fffffffe94ef47e18fbe18c7def7bda53bded3ffffffffffff"),
                (x"fffffffe94ef47e18fbe18c7def7bda53bded3ffffffffffff"),
                (x"ffffffffbdf7463f7bc3f77bdf7bdef77b4a769fffffffffff"),
                (x"ffffffffbd1f7c3f787eed294a5294efbbded280ffffffffff"),
                (x"fffffffe94f53beef69d4def74d294a53bdef680ffffffffff"),
                (x"fffffffe94f53beef69d4def74d294a53bdef680ffffffffff"),
                (x"ffffffffffea7bda52f7bdef7ba7bdef694a5294003fffffff"),
                (x"ffffffffff65ef7bdef7bdef7ba694a77bdef694003fffffff"),
                (x"ffffffffff026f7bdee9eb197ba694a5014a5294003fffffff"),
                (x"ffffffffffa32f74a7bda2529ba7bded28000014003fffffff"),
                (x"fffffffffffd2f7ef69462537bf694ef694a53b4003fffffff"),
                (x"fffffffffffd2f7ef69462537bf694ef694a53b4003fffffff"),
                (x"fffffffffff82f74a4002def7bd3bda769ded3b4003fffffff"),
                (x"fffffffffff82f7bdc0025ef7bd3dea529ded3b4003fffffff"),
                (x"fffffffffff82f7bdf9c25ef7bd3dee8294a769da53fffffff"),
                (x"fffffffffff82f7bddce25ef7bd3dee82800741da53fffffff"),
                (x"fffffffffff82f7bddce25ef7bd3dee82800741da53fffffff"),
                (x"fffffffffff82f7bdef7bdef7bd3dee828007414a53fffffff"),
                (x"fffffffffff8137bdef7bdef74d3dea000005014a53fffffff"),
                (x"ffffffffffffc09bdef7bdee9633bda500000014003fffffff"),
                (x"fffffffffffffe00018c6318cf32940780000014003fffffff"),
                (x"fffffffffffffe00018c6318cf32940780000014003fffffff"),
                (x"ffffffffffffffff780c318cf324004a7c000014003fffffff"),
                (x"ffffffffffffffe7bfd0294be7a4c64dd3ef0000003fffffff"),
                (x"ffffffffffffffef7a102fbde325294defef0000ffffffffff"),
                (x"ffffffffffffffe7bcb0f0000633debdefef7fffffffffffff"),
                (x"ffffffffffffffe7bcb0f0000633debdefef7fffffffffffff"),
                (x"ffffffffffffffe840a502537ba6f7bdee007fffffffffffff"),
                (x"ffffffffffffffe7bcb005ef7bdef7bdd8007fffffffffffff"),
                (x"fffffffffffffff318c602537ba6f7ba41ffffffffffffffff"),
                (x"fffffffffffffffffe86300006318c003fffffffffffffffff"),
                (x"fffffffffffffffffe86300006318c003fffffffffffffffff"),
                (x"fffffffffffffffffe9d39cfdef7bde83fffffffffffffffff"),
                (x"fffffffffffffffffff43bde7ef7bd07ffffffffffffffffff"),
                (x"ffffffffffffffffffffe9cef3f7bd07ffffffffffffffffff"),
                (x"ffffffffffffffffffff03def7f400ffffffffffffffffffff"),
                (x"ffffffffffffffffffff03def7f400ffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc5f7400ffffffffffffffffffff"),

                -- 6_character_1_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ef7bdef7bded29ffffffffffffffff"),
                (x"ffffffffffffff4a53bef0c7eefbdef77b4a53ffffffffffff"),
                (x"ffffffffffffff4a53bef0c7eefbdef77b4a53ffffffffffff"),
                (x"fffffffffffd3bef7bddf0c63f0fdef769def7b4ffffffffff"),
                (x"ffffffffffa77c318fdef0c6318fdef53b4a77dda53fffffff"),
                (x"ffffffffffa53be18c7eefbc318fdeed29defbb4a53fffffff"),
                (x"ffffffffffa53be18c7eefbc318fdeed29defbb4a53fffffff"),
                (x"fffffffc00ef69df787eefbc3f0fdeed3bef769def69ffffff"),
                (x"fffffffc00a7bb4ef7bef77bee8fbda53bded3bea501ffffff"),
                (x"fffffffc00a77dda529df77beefbbda77b4a03dda501ffffff"),
                (x"fffffffc00ed3beef694ef7bda7694a7680053b4a501ffffff"),
                (x"fffffffc00a7694ef694a529da7694a5294a50140001ffffff"),
                (x"fffffffc00a7694ef694a529da7694a5294a50140001ffffff"),
                (x"ffffffffff077bda5294a5294a5294a5294a0294003fffffff"),
                (x"ffffffffff053bdef7b4ed294a5294a528005280003fffffff"),
                (x"ffffffffff053bdef7b4ed294a5294a5294a52800001ffffff"),
                (x"ffffffffff053deef7d4ef7b4a7694a5294a50140001ffffff"),
                (x"ffffffffff053deef7d4ef7b4a7694a5294a50140001ffffff"),
                (x"ffffffffff077dda53d4ef7b4a7694a5294a52940001ffffff"),
                (x"ffffffffffa77d4ef7ddef7bda77bda5294a5294a501ffffff"),
                (x"ffffffffffa77d4ef7ddef7bda77bded294a5280a501ffffff"),
                (x"fffffffffffd3a0ef7d4f7bdda77deed28005280a501ffffff"),
                (x"fffffffffffd3a0ef7d4f7bdda77deed28005280a501ffffff"),
                (x"fffffffffff53a0a53b4efbdda77dee828005280a501ffffff"),
                (x"fffffffffff028000280a7bd4a53dee828005280003fffffff"),
                (x"fffffffffff241000000a77b4053bda028005009f7bfffffff"),
                (x"ffffffffff67bde31a0505294052940400f78129f7bfffffff"),
                (x"ffffffffff67bde31a0505294052940400f78129f7bfffffff"),
                (x"ffffffffff03180319f028000280007bcc94a53e633fffffff"),
                (x"fffffffffff8000f78cf7c2107bfdef781ef7bc9633fffffff"),
                (x"fffffffffffffffa50c6318c6318c631a8c62520ffffffffff"),
                (x"fffffffffffffffa53bd3bdefef4e73f694a001fffffffffff"),
                (x"fffffffffffffffa53bd3bdefef4e73f694a001fffffffffff"),
                (x"fffffffffffffffa529de9ce7ed294a500007fffffffffffff"),
                (x"fffffffffffffffffc14ef7bd383bde83fffffffffffffffff"),
                (x"ffffffffffffffffffe0a1ce7a000007ffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc3f03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bc3f03ffffffffffffffffffffff"),
                (x"ffffffffffffffffffff07bdde83ffffffffffffffffffffff"),

                -- 6_character_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffd8cef7bded294ef694a53ffffffffffff"),
                (x"fffffffffffffecef7bdefbdef7bdea0fddef694ffffffffff"),
                (x"fffffffffffffecef7bdefbdef7bdea0fddef694ffffffffff"),
                (x"ffffffffffffe9def694ef7bde8c63f747ef0fbda53fffffff"),
                (x"fffffffffffd3b4ef7bef7bdeef7de1fbc318fbeef7fffffff"),
                (x"ffffffffff0529def7dda5294a53bdf0fc31fba3ef7fffffff"),
                (x"ffffffffff0529def7dda5294a53bdf0fc31fba3ef7fffffff"),
                (x"ffffffffff053bdef694a5289bdd29ed3bef769ea53fffffff"),
                (x"fffffffc00a5294a53bdea537bdef7bde9def53dffffffffff"),
                (x"fffffffc00a53bdef7b4a2537bdef7bdef7bdeecffffffffff"),
                (x"fffffffc00a529400294a2537bb3bd4def7bdd20ffffffffff"),
                (x"fffffffc00a7680a529dea5374a694ef537bdd94ffffffffff"),
                (x"fffffffc00a7680a529dea5374a694ef537bdd94ffffffffff"),
                (x"fffffffc00ed3b4a53bda77b7ba58ca53b7bde9fffffffffff"),
                (x"ffffff8294ed3b4003b4ed297bdca500137bdc1fffffffffff"),
                (x"ffffff83bda77b400294f5297bdc84002f7bdc1fffffffffff"),
                (x"ffffff83bda76800001df5297bdc84e72f7bdc1fffffffffff"),
                (x"ffffff83bda76800001df5297bdc84e72f7bdc1fffffffffff"),
                (x"ffffff83bda76800001df77b7bdc8473af7bdc1fffffffffff"),
                (x"fffff053bda768000014f77b7bdef7bdef7bdc1fffffffffff"),
                (x"fffff05294ed00000014efbccbdef7bdef7ba41fffffffffff"),
                (x"fffff05000ed00000280a77ac4def7bdee9483ffffffffffff"),
                (x"fffff05000ed00000280a77ac4def7bdee9483ffffffffffff"),
                (x"ffffffd000a0000003c90528c6318c6300007fffffffffffff"),
                (x"ffffff8000a0000002f748009f18c6303dffffffffffffffff"),
                (x"fffffffc00003e0f7af74a52934210879e007fffffffffffff"),
                (x"ffffffffff003e0f7937ba529f3e10878c007fffffffffffff"),
                (x"ffffffffff003e0f7937ba529f3e10878c007fffffffffffff"),
                (x"fffffffffffffe0318d7bdefef0000019fef7fffffffffffff"),
                (x"fffffffffffffe031bc9bdee965ef7b81fef7fffffffffffff"),
                (x"fffffffffffffe0f78c04def74def7b80def7fffffffffffff"),
                (x"ffffffffffffffd003de025374a6f76741ffffffffffffffff"),
                (x"ffffffffffffffd003de025374a6f76741ffffffffffffffff"),
                (x"ffffffffffffffdef4e7e800c60000077fffffffffffffffff"),
                (x"fffffffffffffe0ef4ef3f7bd077bdefffffffffffffffffff"),
                (x"fffffffffffffe0ef7a7ef7bd074e73f7fffffffffffffffff"),
                (x"fffffffffffffff000ef3f7a0003bdf7bfffffffffffffffff"),
                (x"fffffffffffffff000ef3f7a0003bdf7bfffffffffffffffff"),
                (x"fffffffffffffff003be2fbc0fffffffffffffffffffffffff"),

                -- 6_character_1_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ef7bdef7bded29ffffffffffffffff"),
                (x"ffffffffffffff4a53bdf0c7eefbdef77b4a53ffffffffffff"),
                (x"ffffffffffffff4a53bdf0c7eefbdef77b4a53ffffffffffff"),
                (x"fffffffffffd3beef69ee8c63f0fdeef69def7b4ffffffffff"),
                (x"ffffffffffa77c3f7bb4f77a318fdeed3b4a77dda53fffffff"),
                (x"ffffffffffa53be18fddf77be1fbbda529defbb4a53fffffff"),
                (x"ffffffffffa53be18fddf77be1fbbda529defbb4a53fffffff"),
                (x"fffffffc00ef69d18fb4a77bdf77bda53bef769def41ffffff"),
                (x"fffffffc00a7bb4ef5374d29def6944dd34a53bea501ffffff"),
                (x"fffffffc00a77d4bdef7bdee9ea6f7bdef7bd3dda501ffffff"),
                (x"fffffffc00a03b4bdef7bdef7bdef7bdef7bd3b4a501ffffff"),
                (x"fffffffc00a7414633a9bdef7bdef7ba7ac6529da501ffffff"),
                (x"fffffffc00a7414633a9bdef7bdef7ba7ac6529da501ffffff"),
                (x"ffffffffffa76894a69dea537bdd29ef6894a41da53fffffff"),
                (x"ffffffffff077dd4a594a77b7bdfbda51894d3b4003fffffff"),
                (x"ffffffffff077d4bdca002537bdd29000b7bd3d4003fffffff"),
                (x"ffffffffff053d4bdc8005ef7bdef700097bd3d4003fffffff"),
                (x"ffffffffff053d4bdc8005ef7bdef700097bd3d4003fffffff"),
                (x"ffffffffffa53a0bdc9ce5ef7bdef7e7097bd3d4a53fffffff"),
                (x"ffffffffffa03a0bdc8e75ef7bdef773897b83a0ef69ffffff"),
                (x"ffffffffffa03a04a6f7bdef7bdef7bdee9483a0ef69ffffff"),
                (x"ffffffffff3028063137bdef7bdef7bdd2c60280f7ba0fffff"),
                (x"ffffffffff3028063137bdef7bdef7bdd2c60280f7ba0fffff"),
                (x"fffffffcc64a6807bc0c4a537bdd294b006302894a7c0fffff"),
                (x"fffffff9294a520840c53318c6318c340cf781294a53efffff"),
                (x"fffffff9294a5267bcc5294be4f8a52c0c6341294a53efffff"),
                (x"ffffffb1294a52031a05294aff3ca529606301294a7dffffff"),
                (x"ffffffb1294a52031a05294aff3ca529606301294a7dffffff"),
                (x"ffffffb1294a58031a05294a5294a529400032f74a59ffffff"),
                (x"ffffffb2f7ba41f319e5294a5294a52bd97bdee94a59ffffff"),
                (x"ffffffb129bb01fef7c6318c6318c637997bdd2c6301ffffff"),
                (x"ffffff81294b3ffef4e77bdef79ce73f4094dd80003fffffff"),
                (x"ffffff81294b3ffef4e77bdef79ce73f4094dd80003fffffff"),
                (x"fffffffc00003ffef7a77bde7ef7bdef7a00001fffffffffff"),
                (x"ffffffffffffffffffa73bde7383bdef7bffffffffffffffff"),
                (x"fffffffffffffffffffd7bdef383bdef7fffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7bde800007ffffffffffffffffff"),
                (x"ffffffffffffffffffe0ef7bde800007ffffffffffffffffff"),
                (x"ffffffffffffffffffffef7beeffffffffffffffffffffffff"),

                -- 6_character_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffe94a53bda529def7bda53fffffffffffffffff"),
                (x"ffffffffffa53bdf7874f7bdef7bbdef7b4a7fffffffffffff"),
                (x"ffffffffffa53bdf7874f7bdef7bbdef7b4a7fffffffffffff"),
                (x"fffffffe94ef47e18fbe18c7def7bda53bded3ffffffffffff"),
                (x"ffffffffbdf7463f7bc3f77bdf7bdef77b4a769fffffffffff"),
                (x"ffffffffbd1f7c3f787eed294a5294efbbded280ffffffffff"),
                (x"ffffffffbd1f7c3f787eed294a5294efbbded280ffffffffff"),
                (x"fffffffe94f53beef69d4def74d294a53bdef680ffffffffff"),
                (x"ffffffffffea7bda52f7bdef7ba7bdef694a5294003fffffff"),
                (x"ffffffffff65ef7bdef7bdef7ba694a77bdef694003fffffff"),
                (x"ffffffffff026f7bdee9eb197ba694a5014a5294003fffffff"),
                (x"ffffffffffa32f74a7bda2529ba7bded280053b4003fffffff"),
                (x"ffffffffffa32f74a7bda2529ba7bded280053b4003fffffff"),
                (x"fffffffffffd2f7ef69462537bf694ef694a769d003fffffff"),
                (x"fffffffffff82f74a4002def7bd3bda7414a769da501ffffff"),
                (x"fffffffffff82f7bdc0025ef7bd3dea5014a77b4ef41ffffff"),
                (x"fffffffffff82f7bdf9c25ef7bd3dee8000053b4ef41ffffff"),
                (x"fffffffffff82f7bdf9c25ef7bd3dee8000053b4ef41ffffff"),
                (x"fffffffffff82f7bddce25ef7bf7dee8000053b4ef41ffffff"),
                (x"fffffffffff82f7bdef7bdef7bf7dea0000053b4ef680fffff"),
                (x"fffffffffff8137bdef7bdef767bbda00000029da5280fffff"),
                (x"ffffffffffffc09bdef7bdee967694050000029d00280fffff"),
                (x"ffffffffffffc09bdef7bdee967694050000029d00280fffff"),
                (x"fffffffffffffe00018c6318c650004f800000140029ffffff"),
                (x"ffffffffffffffff7806318de48129ba400000140001ffffff"),
                (x"fffffffffffffe07be1087bc64a6f7ba7c007c00003fffffff"),
                (x"fffffffffffffe031a10f3dfe4a6f7ba7c007c00ffffffffff"),
                (x"fffffffffffffe031a10f3dfe4a6f7ba7c007c00ffffffffff"),
                (x"ffffffffffffffe7bcc00001ef5ef7b98c007fffffffffffff"),
                (x"ffffffffffffffe7bc17bdeec4def74f8c007fffffffffffff"),
                (x"ffffffffffffffe31817bdee9bdd2901bc007fffffffffffff"),
                (x"fffffffffffffff003acba529ba400f781deffffffffffffff"),
                (x"fffffffffffffff003acba529ba400f781deffffffffffffff"),
                (x"ffffffffffffffffffa00000c603bd39fbdeffffffffffffff"),
                (x"fffffffffffffffffffdef7a0ef4e779fa007fffffffffffff"),
                (x"ffffffffffffffffffa73f7a0ef7bd3f7a007fffffffffffff"),
                (x"ffffffffffffffffffdee8000074e779c1ffffffffffffffff"),
                (x"ffffffffffffffffffdee8000074e779c1ffffffffffffffff"),
                (x"fffffffffffffffffffffffff078a5f741ffffffffffffffff"),

                -- 6_character_2_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ef7bdef7bded29ffffffffffffffff"),
                (x"ffffffffffffff4a53bef0c7eefbdef77b4a53ffffffffffff"),
                (x"ffffffffffffff4a53bef0c7eefbdef77b4a53ffffffffffff"),
                (x"fffffffffffd3bef7bddf0c63f0fdef769def7b4ffffffffff"),
                (x"ffffffffffa77c318fdef0c6318fdef53b4a77dda53fffffff"),
                (x"ffffffffffa53be18c7eefbc318fdeed29defbb4a53fffffff"),
                (x"ffffffffffa53be18c7eefbc318fdeed29defbb4a53fffffff"),
                (x"fffffffc00ef69df787eefbc3f0fdeed3bef769def69ffffff"),
                (x"fffffffc00a7bb4ef7bef77bee8fbda53bded3bea501ffffff"),
                (x"fffffffc00a77dda529df77beefbbda77b4a03dda501ffffff"),
                (x"fffffffc00ed3beef694ef7bda7694a7680053b4a501ffffff"),
                (x"fffffffc00a7694ef694a529da7694a5294a50140001ffffff"),
                (x"fffffffc00a7694ef694a529da7694a5294a50140001ffffff"),
                (x"ffffffffff077bda5294a5294a5294a5294a0294003fffffff"),
                (x"ffffffffff077bdef694ed294a5294a528005280003fffffff"),
                (x"ffffffffffa77bdef694ef7bda5294a5294a5000003fffffff"),
                (x"ffffffffffa77bdef69def7bda5294a5294a5280003fffffff"),
                (x"ffffffffffa77bdef69def7bda5294a5294a5280003fffffff"),
                (x"ffffffffffa77beef69def7bda7694a7694a5280003fffffff"),
                (x"fffffffe94f769eef69def7bda7694a7694a0280003fffffff"),
                (x"fffffffe94f53beef69de801def694a7694a0280ffffffffff"),
                (x"ffffffffdeed3dda53bee801df7694ef68005280ffffffffff"),
                (x"ffffffffdeed3dda53bee801df7694ef68005280ffffffffff"),
                (x"ffffffffbd053d4a53dea001df7694ef68005280f7bfffffff"),
                (x"fffffffe9400280a53dda0014f5000ed28005009f7bfffffff"),
                (x"fffffffffff2400a53dd00014ed000ed014a5009f7bfffffff"),
                (x"fffffffffff2529003b400014a0000a0000003de633fffffff"),
                (x"fffffffffff2529003b400014a0000a0000003de633fffffff"),
                (x"ffffffffff679294a4007c200014a5001e63018c003fffffff"),
                (x"ffffffffff627def781ef7bcf7c2107bcdef0000ffffffffff"),
                (x"fffffffffff81296329def7bde98c6318d4a7fffffffffffff"),
                (x"ffffffffffffc00a529d39cfdebdef3f7b4a7fffffffffffff"),
                (x"ffffffffffffc00a529d39cfdebdef3f7b4a7fffffffffffff"),
                (x"fffffffffffffff00014a5294e9ce7ef694a7fffffffffffff"),
                (x"ffffffffffffffffffe0ef7a03f7bded01ffffffffffffffff"),
                (x"ffffffffffffffffffff00000a1ce7a03fffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f0fde07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0f0fde07ffffffffffffffffff"),
                (x"fffffffffffffffffffffffe0ef7de07ffffffffffffffffff"),

                -- 6_character_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ef7bded294ef694a53ffffffffffff"),
                (x"ffffffffffffff4ef7bdefbdef7bdea0fddef694ffffffffff"),
                (x"ffffffffffffff4ef7bdefbdef7bdea0fddef694ffffffffff"),
                (x"ffffffffffffe9def694ef7bde8c63f747ef0fbda53fffffff"),
                (x"fffffffffffd3b4ef7bef7bdeef7de1fbc318fbeef7fffffff"),
                (x"ffffffffff0529def7dda5294a53bdf0fc31fba3ef7fffffff"),
                (x"ffffffffff0529def7dda5294a53bdf0fc31fba3ef7fffffff"),
                (x"ffffffffff053bdef694a5289bdd29ed3bef769ea53fffffff"),
                (x"fffffffc00a5294a53bdea537bdef7bde9def53dffffffffff"),
                (x"fffffffc00a53bdef7b4a2537bdef7bdef7bdeecffffffffff"),
                (x"fffffffc00a5294a5294a2537bb3bd4def7bdd20ffffffffff"),
                (x"fffffffc00053b4a501dea5374a694ef537bdd94ffffffffff"),
                (x"fffffffc00053b4a501dea5374a694ef537bdd94ffffffffff"),
                (x"fffffffc00053b4a53bda77b7ba58ca53b7bde9fffffffffff"),
                (x"fffffffc00a53b4a53b4ed297bdca500137bdc1fffffffffff"),
                (x"fffffffc00a769da5294f5297bdc84002f7bdc1fffffffffff"),
                (x"fffffffe94a769da501df5297bdc84e72f7bdc1fffffffffff"),
                (x"fffffffe94a769da501df5297bdc84e72f7bdc1fffffffffff"),
                (x"fffffffe94a76940001df5297bdc8473af7bdc1fffffffffff"),
                (x"fffffffe94a74140001df5297bdef7bdef7bdc1fffffffffff"),
                (x"fffffffe94a740000014f5289bdef7bdef7ba41fffffffffff"),
                (x"fffffffc00a740000294eb18c4def7bdee9483ffffffffffff"),
                (x"fffffffc00a740000294eb18c4def7bdee9483ffffffffffff"),
                (x"fffffffc00a740000120a319e6318c6300007fffffffffffff"),
                (x"ffffffffff050004a6e9018cf818c6483dffffffffffffffff"),
                (x"ffffffffff0501ebdee94bdfe29610f41fef7fffffffffffff"),
                (x"fffffffffff8006bdee94bdef84210879ec67fffffffffffff"),
                (x"fffffffffff8006bdee94bdef84210879ec67fffffffffffff"),
                (x"ffffffffffffc09bdef74fbc68421083fc94b3ffffffffffff"),
                (x"ffffffffffffc1e4a6f7480008421083fc9483ffffffffffff"),
                (x"fffffffffffffe04a6f7bdee9f3def7f80007fffffffffffff"),
                (x"fffffffffffffe063137bdef7018c63181ffffffffffffffff"),
                (x"fffffffffffffe063137bdef7018c63181ffffffffffffffff"),
                (x"fffffffffffffff0000c4dee903def3f7fffffffffffffffff"),
                (x"fffffffffffffff003bd00000e9fbdef7fffffffffffffffff"),
                (x"fffffffffffffffef7bd00000e9def79ffffffffffffffffff"),
                (x"fffffffffffffff0001de8000074e7ef41ffffffffffffffff"),
                (x"fffffffffffffff0001de8000074e7ef41ffffffffffffffff"),
                (x"fffffffffffffffffffffffff077de2f81ffffffffffffffff"),

                -- 6_character_2_2
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffe94ef7bdef7bded29ffffffffffffffff"),
                (x"ffffffffffffff4a53bdf0c7eefbdef77b4a53ffffffffffff"),
                (x"ffffffffffffff4a53bdf0c7eefbdef77b4a53ffffffffffff"),
                (x"fffffffffffd3beef69ee8c63f0fdeef69def7b4ffffffffff"),
                (x"ffffffffffa77c3f7bb4f77a318fdeed3b4a77dda53fffffff"),
                (x"ffffffffffa53be18fddf77be1fbbda529defbb4a53fffffff"),
                (x"ffffffffffa53be18fddf77be1fbbda529defbb4a53fffffff"),
                (x"fffffffc00ef69d18fb4a77bdf77bda53bef769def41ffffff"),
                (x"fffffffc00a7bb4ef5374d29def6944dd34a53bea501ffffff"),
                (x"fffffffc00a77d4bdef7bdee9ea6f7bdef7bd3dda501ffffff"),
                (x"fffffffc00a03b4bdef7bdef7bdef7bdef7bd3b4a501ffffff"),
                (x"fffffffc00a7414633a9bdef7bdef7ba7ac6529da501ffffff"),
                (x"fffffffc00a7414633a9bdef7bdef7ba7ac6529da501ffffff"),
                (x"ffffffffffa76894a69dea537bdd29ef6894a41da53fffffff"),
                (x"ffffffffff077dd4a594a77b7bdfbda51894d3b4003fffffff"),
                (x"ffffffffff077d4bdca002537bdd29000b7bd3d4003fffffff"),
                (x"ffffffffff053d4bdc8005ef7bdef700097bd3d4003fffffff"),
                (x"ffffffffff053d4bdc8005ef7bdef700097bd3d4003fffffff"),
                (x"fffffffe94a53a0bdc9ce5ef7bdef7e7097bd3d4a53fffffff"),
                (x"fffffffe94e83a0bdc8e75ef7bdef773897b83a0a53fffffff"),
                (x"fffffffe94e83a04a6f7bdef7bdef7bdee9483a0a53fffffff"),
                (x"ffffffd3bdf028063137bdef7bdef7bdd2c6028031bfffffff"),
                (x"ffffffd3bdf028063137bdef7bdef7bdd2c6028031bfffffff"),
                (x"fffffffbde4a6803180c4a537bdd294b00f782894a4dffffff"),
                (x"fffffff9294a5207bcd03318c6318c314d0801294a53efffff"),
                (x"fffffff9294a529318d0294be4f8a52c0cf799294a53efffff"),
                (x"fffffff9294a52031a05294aff3ca529606301296312cfffff"),
                (x"fffffff9294a52031a05294aff3ca529606301296312cfffff"),
                (x"fffffffd8c4deec00005294a5294a5296063018c4a52cfffff"),
                (x"fffffffd8c4a6f7bdd8f294a5294a5295e637c09bdeecfffff"),
                (x"fffffffc0063137bdd9e318c6318c67fbddefc0cbdd2cfffff"),
                (x"ffffffffff001974a41d39ce77bdef79cfdeffec4a520fffff"),
                (x"ffffffffff001974a41d39ce77bdef79cfdeffec4a520fffff"),
                (x"ffffffffffffc00003bdef7bde9def79fbdeffe00001ffffff"),
                (x"ffffffffffffffffffbdef7a039def39fbffffffffffffffff"),
                (x"fffffffffffffffffffdef7a03bdef7f7fffffffffffffffff"),
                (x"ffffffffffffffffffff00000ef7bde83fffffffffffffffff"),
                (x"ffffffffffffffffffff00000ef7bde83fffffffffffffffff"),
                (x"fffffffffffffffffffffffffefbbdefffffffffffffffffff"),

                -- 6_character_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffe94a53bda529def7bda53fffffffffffffffff"),
                (x"ffffffffffa53bdf7874f7bdef7bbdef7b4a7fffffffffffff"),
                (x"ffffffffffa53bdf7874f7bdef7bbdef7b4a7fffffffffffff"),
                (x"fffffffe94ef47e18fbe18c7def7bda53bded3ffffffffffff"),
                (x"ffffffffbdf7463f7bc3f77bdf7bdef77b4a769fffffffffff"),
                (x"ffffffffbd1f7c3f787eed294a5294efbbded280ffffffffff"),
                (x"ffffffffbd1f7c3f787eed294a5294efbbded280ffffffffff"),
                (x"fffffffe94f53beef69d4def74d294a53bdef680ffffffffff"),
                (x"ffffffffffea7bda52f7bdef7ba7bdef694a5294003fffffff"),
                (x"ffffffffff65ef7bdef7bdef7ba694a77bdef694003fffffff"),
                (x"ffffffffff026f7bdee9eb197ba694a5294a5294003fffffff"),
                (x"ffffffffffa32f74a7bda2529ba7bde8294a7680003fffffff"),
                (x"ffffffffffa32f74a7bda2529ba7bde8294a7680003fffffff"),
                (x"fffffffffffd2f7ef69462537bf694ef694a7680003fffffff"),
                (x"fffffffffff82f74a4002def7bd3bda7694a7694003fffffff"),
                (x"fffffffffff82f7bdc0025ef7bd3dea529ded3b4003fffffff"),
                (x"fffffffffff82f7bdf9c25ef7bd3dee829ded3b4a53fffffff"),
                (x"fffffffffff82f7bdf9c25ef7bd3dee829ded3b4a53fffffff"),
                (x"fffffffffff82f7bddce25ef7bd3dee8014a53b4a53fffffff"),
                (x"fffffffffff82f7bdef7bdef7bd3dee8014a03b4a53fffffff"),
                (x"fffffffffff8137bdef7bdef74d3dea0000003b4a53fffffff"),
                (x"ffffffffffffc09bdef7bdee9633bda5000003b4003fffffff"),
                (x"ffffffffffffc09bdef7bdee9633bda5000003b4003fffffff"),
                (x"fffffffffffffe00018c6318cf329402400003b4003fffffff"),
                (x"ffffffffffffffff7809318d0798004dee000280ffffffffff"),
                (x"ffffffffffffffe7be1e814a5f3d294defef0280ffffffffff"),
                (x"fffffffffffffec7bfcf814b07bd294dee94801fffffffffff"),
                (x"fffffffffffffec7bfcf814b07bd294dee94801fffffffffff"),
                (x"ffffffffffffd89f79f08421037a104dee9483ffffffffffff"),
                (x"ffffffffffffc09f79f08421000129bdd3ef03ffffffffffff"),
                (x"fffffffffffffe0003cf7bdfe4def7bdd2007fffffffffffff"),
                (x"fffffffffffffff000c6318c0bdef7ba58007fffffffffffff"),
                (x"fffffffffffffff000c6318c0bdef7ba58007fffffffffffff"),
                (x"ffffffffffffffffffa77bde04dd296001ffffffffffffffff"),
                (x"ffffffffffffffffffbde9cfd00000ef41ffffffffffffffff"),
                (x"fffffffffffffffffcef79cfd00000ef7bffffffffffffffff"),
                (x"fffffffffffffff003bd3f7a0003bde801ffffffffffffffff"),
                (x"fffffffffffffff003bd3f7a0003bde801ffffffffffffffff"),
                (x"fffffffffffffff003c5f77a0fffffffffffffffffffffffff")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 3359 := 0;
    signal out_color_reg : std_logic_vector(199 downto 0) := (others => '0');
begin
    process(in_sprite_id, in_sprite_row, in_sprite_col, in_sprite_state, in_sprite_direction)
    begin
        real_row <= 0;
        case in_sprite_id is
            when 0 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= in_sprite_row;
                            when D_LEFT => real_row <= 40 + in_sprite_row;
                            when D_DOWN => real_row <= 80 + in_sprite_row;
                            when D_RIGHT => real_row <= 120 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 160 + in_sprite_row;
                            when D_LEFT => real_row <= 200 + in_sprite_row;
                            when D_DOWN => real_row <= 240 + in_sprite_row;
                            when D_RIGHT => real_row <= 280 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 320 + in_sprite_row;
                            when D_LEFT => real_row <= 360 + in_sprite_row;
                            when D_DOWN => real_row <= 400 + in_sprite_row;
                            when D_RIGHT => real_row <= 440 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 1 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 480 + in_sprite_row;
                            when D_LEFT => real_row <= 520 + in_sprite_row;
                            when D_DOWN => real_row <= 560 + in_sprite_row;
                            when D_RIGHT => real_row <= 600 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 640 + in_sprite_row;
                            when D_LEFT => real_row <= 680 + in_sprite_row;
                            when D_DOWN => real_row <= 720 + in_sprite_row;
                            when D_RIGHT => real_row <= 760 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 800 + in_sprite_row;
                            when D_LEFT => real_row <= 840 + in_sprite_row;
                            when D_DOWN => real_row <= 880 + in_sprite_row;
                            when D_RIGHT => real_row <= 920 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 2 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 960 + in_sprite_row;
                            when D_LEFT => real_row <= 1000 + in_sprite_row;
                            when D_DOWN => real_row <= 1040 + in_sprite_row;
                            when D_RIGHT => real_row <= 1080 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1120 + in_sprite_row;
                            when D_LEFT => real_row <= 1160 + in_sprite_row;
                            when D_DOWN => real_row <= 1200 + in_sprite_row;
                            when D_RIGHT => real_row <= 1240 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1280 + in_sprite_row;
                            when D_LEFT => real_row <= 1320 + in_sprite_row;
                            when D_DOWN => real_row <= 1360 + in_sprite_row;
                            when D_RIGHT => real_row <= 1400 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 3 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1440 + in_sprite_row;
                            when D_LEFT => real_row <= 1480 + in_sprite_row;
                            when D_DOWN => real_row <= 1520 + in_sprite_row;
                            when D_RIGHT => real_row <= 1560 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1600 + in_sprite_row;
                            when D_LEFT => real_row <= 1640 + in_sprite_row;
                            when D_DOWN => real_row <= 1680 + in_sprite_row;
                            when D_RIGHT => real_row <= 1720 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1760 + in_sprite_row;
                            when D_LEFT => real_row <= 1800 + in_sprite_row;
                            when D_DOWN => real_row <= 1840 + in_sprite_row;
                            when D_RIGHT => real_row <= 1880 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 4 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1920 + in_sprite_row;
                            when D_LEFT => real_row <= 1960 + in_sprite_row;
                            when D_DOWN => real_row <= 2000 + in_sprite_row;
                            when D_RIGHT => real_row <= 2040 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2080 + in_sprite_row;
                            when D_LEFT => real_row <= 2120 + in_sprite_row;
                            when D_DOWN => real_row <= 2160 + in_sprite_row;
                            when D_RIGHT => real_row <= 2200 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2240 + in_sprite_row;
                            when D_LEFT => real_row <= 2280 + in_sprite_row;
                            when D_DOWN => real_row <= 2320 + in_sprite_row;
                            when D_RIGHT => real_row <= 2360 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 5 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2400 + in_sprite_row;
                            when D_LEFT => real_row <= 2440 + in_sprite_row;
                            when D_DOWN => real_row <= 2480 + in_sprite_row;
                            when D_RIGHT => real_row <= 2520 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2560 + in_sprite_row;
                            when D_LEFT => real_row <= 2600 + in_sprite_row;
                            when D_DOWN => real_row <= 2640 + in_sprite_row;
                            when D_RIGHT => real_row <= 2680 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2720 + in_sprite_row;
                            when D_LEFT => real_row <= 2760 + in_sprite_row;
                            when D_DOWN => real_row <= 2800 + in_sprite_row;
                            when D_RIGHT => real_row <= 2840 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 6 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 2880 + in_sprite_row;
                            when D_LEFT => real_row <= 2920 + in_sprite_row;
                            when D_DOWN => real_row <= 2960 + in_sprite_row;
                            when D_RIGHT => real_row <= 3000 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 3040 + in_sprite_row;
                            when D_LEFT => real_row <= 3080 + in_sprite_row;
                            when D_DOWN => real_row <= 3120 + in_sprite_row;
                            when D_RIGHT => real_row <= 3160 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 3200 + in_sprite_row;
                            when D_LEFT => real_row <= 3240 + in_sprite_row;
                            when D_DOWN => real_row <= 3280 + in_sprite_row;
                            when D_RIGHT => real_row <= 3320 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= rom(real_row);
        end if;
    end process;
    out_color <= out_color_reg(((in_sprite_col + 1) * 5) - 1 downto (in_sprite_col * 5));
end behavioral;
