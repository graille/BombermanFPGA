library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.PROJECT_PARAMS_PKG.all;
use work.PROJECT_TYPES_PKG.all;
use work.PROJECT_DIRECTION_PKG.all;

entity ressources_sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_id : in block_category_type;
        in_sprite_state : in state_type;
        in_sprite_direction : in direction_type;

        in_sprite_row : in integer range 0 to 39;
        in_sprite_col : in integer range 0 to 39;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end ressources_sprite_rom;

architecture behavioral of ressources_sprite_rom is
    subtype word_t is std_logic_vector(0 to 199);
    type memory_t is array(0 to 1719) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- 0_empty
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 1_unbreakable
                (x"ef7af784210842108421084210842108421084210842118def"),
                (x"ef7af784210842108421084210842108421084210842118def"),
                (x"ef7af784210842108421084210842108421084210842118def"),
                (x"ef7af790840842108421084210842108421084210908418def"),
                (x"ef7af790840842108421084210842108421084210908418def"),
                (x"ef7af784210848421084210842108421084210210842118def"),
                (x"ef7af784210848421084210842108421084210210842118def"),
                (x"ef7af784210848421084210842108421084210210842118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784212108421084210842108421084210842042118def"),
                (x"ef7af784210848421084210842108421084210210842118def"),
                (x"ef7af784210848421084210842108421084210210842118def"),
                (x"ef7af790840842108421084210842108421084210908418def"),
                (x"ef7af790840842108421084210842108421084210908418def"),
                (x"ef7af790840842108421084210842108421084210908418def"),
                (x"ef7af78c6318c6318c6318c6318c6318c6318c6318c6318def"),
                (x"ef7af78c6318c6318c6318c6318c6318c6318c6318c6318def"),
                (x"ef7bef3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef"),
                (x"ef7bef3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef"),
                (x"ef7bef3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef"),
                (x"ef7bdefbdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde"),
                (x"ef7bdefbdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde"),
                (x"ef7bdefbdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde"),
                (x"ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7de"),
                (x"ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7de"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce739c"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce739c"),

                -- 2_unbreakable
                (x"e739def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e739def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e739def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e738f790842108421084210842108421084210842108418fbd"),
                (x"e738f790842108421084210842108421084210842108418fbd"),
                (x"e739ef0c6308421084210842108421084210842108c637bfbd"),
                (x"e739ef0c6308421084210842108421084210842108c637bfbd"),
                (x"e739ef0c6308421084210842108421084210842108c637bfbd"),
                (x"e739ef3def085ef7bdef7bdef7bdef7bdef7bc2108c637bfbd"),
                (x"e739ef3def085ef7bdef7bdef7bdef7bdef7bc2108c637bfbd"),
                (x"e739ef3def08463190842106318c64210847bc2108c637bfbd"),
                (x"e739ef3def08463190842106318c64210847bc2108c637bfbd"),
                (x"e739ef3def08463190842106318c64210847bc2108c637bfbd"),
                (x"e739ef3def084631bdef2106318c6f790847bc2108c637bfbd"),
                (x"e739ef3def084631bdef2106318c6f790847bc2108c637bfbd"),
                (x"e739ef3def084631bdef2106318c6f790847bc2108c637bfbd"),
                (x"e739ef3def0846318c6318c6318c6318c637bc2108c637bfbd"),
                (x"e739ef3def0846318c6318c6318c6318c637bc2108c637bfbd"),
                (x"e739ef3def08463190842106318c64210847bc2108c637bfbd"),
                (x"e739ef3def08463190842106318c64210847bc2108c637bfbd"),
                (x"e739ef3def084631bdef2106318c6f790847bc2108c637bfbd"),
                (x"e739ef3def084631bdef2106318c6f790847bc2108c637bfbd"),
                (x"e739ef3def084631bdef2106318c6f790847bc2108c637bfbd"),
                (x"e739ef3def0846318c6318c6318c6318c637bc2108c637bfbd"),
                (x"e739ef3def0846318c6318c6318c6318c637bc2108c637bfbd"),
                (x"e739ef3def08421084210842108421084210842108c637bfbd"),
                (x"e739ef3def08421084210842108421084210842108c637bfbd"),
                (x"e739ef3def08421084210842108421084210842108c637bfbd"),
                (x"e739ef3def18c6318c6318c6318c6318c6318c6318c637bfbd"),
                (x"e739ef3def18c6318c6318c6318c6318c6318c6318c637bfbd"),
                (x"e739ef3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bfbd"),
                (x"e739ef3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bfbd"),
                (x"e739ef3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bfbd"),
                (x"e739ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde7bfbd"),
                (x"e739ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde7bfbd"),
                (x"e739ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde7bfbd"),
                (x"e739def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e739def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce73bd"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce73bd"),

                -- 3_breakable
                (x"318c42108421084210842108421084218c639c6318c6318c63"),
                (x"318c42108421084210842108421084218c639c6318c6318c63"),
                (x"318c42108421084210842108421084218c639c6318c6318c63"),
                (x"39ce4210842108421084210842108421ce739c6318c6318c63"),
                (x"39ce4210842108421084210842108421ce739c6318c6318c63"),
                (x"39ce4210842108421084210842108421ce739c6318c6318c63"),
                (x"39ce4210842108421084210842108421ce739c6318c6318c63"),
                (x"39ce4210842108421084210842108421ce739c6318c6318c63"),
                (x"39ce42108421084210842108421084218c639c6318c6318c63"),
                (x"39ce42108421084210842108421084218c639c6318c6318c63"),
                (x"39ce5294a5294a5294a5294a5294a5298c639ce739ce739ce7"),
                (x"39ce5294a5294a5294a5294a5294a5298c639ce739ce739ce7"),
                (x"39ce5294a5294a5294a5294a5294a5298c639ce739ce739ce7"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"294a5294a5318a52908421084210842108421084218c618ca5"),
                (x"294a5294a5318a52908421084210842108421084218c618ca5"),
                (x"294a5294a5318a5290842108421084210842108421ce718ca5"),
                (x"294a5294a5318a5290842108421084210842108421ce718ca5"),
                (x"18c6318c6339ca5290842108421084210842108421ce718c63"),
                (x"18c6318c6339ca5290842108421084210842108421ce718c63"),
                (x"18c6318c6339ca5290842108421084210842108421ce718c63"),
                (x"18c6318c63318a5294a5294a5294a5294a5294a529ce718c63"),
                (x"18c6318c63318a5294a5294a5294a5294a5294a529ce718c63"),
                (x"39ce6318c6318c631ce7318c6318c6318c6318c631ce739ce7"),
                (x"39ce6318c6318c631ce7318c6318c6318c6318c631ce739ce7"),
                (x"39ce6318c6318c631ce7318c6318c6318c6318c631ce739ce7"),
                (x"2108421084210842108439c6318c6318c6318cc63108421084"),
                (x"2108421084210842108439c6318c6318c6318cc63108421084"),
                (x"2108421084210842108439c6318c6318c6318cc63108421084"),
                (x"2108421084210842108439c6318c6318c6318cc63108421084"),
                (x"2108421084210842108439c6318c6318c6318cc63108421084"),
                (x"294a5294a5294a5294a539c6318c6318c6318cc6314a5294a5"),
                (x"294a5294a5294a5294a539c6318c6318c6318cc6314a5294a5"),
                (x"294a5294a5294a5294a539c6318c6318c6318cc6314a5294a5"),
                (x"39ce739ce739ce739ce739ce739ce739ce739cc631ce739ce7"),
                (x"39ce739ce739ce739ce739ce739ce739ce739cc631ce739ce7"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),

                -- 4_bomb_0
                (x"fffffffffffffffffffffffffffffffffffffffffa108fffff"),
                (x"fffffffffffffffffffffffffffffffffffffffffa108fffff"),
                (x"fffffffffffffffffffffffffffffffffffffffffa108fffff"),
                (x"ffffffffffffffffffe000000000000000007fe004e73423ff"),
                (x"ffffffffffffffffffe000000000000000007fe004e73423ff"),
                (x"ffffffffffffc000001ce739ce739ce73fff801ff8000fffff"),
                (x"ffffffffffffc000001ce739ce739ce73fff801ff8000fffff"),
                (x"ffffffffffffc000001ce739ce739ce73fff801ff8000fffff"),
                (x"ffffffffff000c6318c1098dce739c0840007fe000000fffff"),
                (x"ffffffffff000c6318c1098dce739c0840007fe000000fffff"),
                (x"ffffff800031a318c631898c631b9c084000001ce739c003ff"),
                (x"ffffff800031a318c631898c631b9c084000001ce739c003ff"),
                (x"ffffff80008c4210842b5c62631b9cfffffff39ce739c003ff"),
                (x"ffffff80008c4210842b5c62631b9cfffffff39ce739c003ff"),
                (x"ffffff80008c4210842b5c62631b9cfffffff39ce739c003ff"),
                (x"fffe0018c68c4210842b5c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c68c4210842b5c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c68c56b5ad6b5c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c68c56b5ad6b5c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c68c6318c6318c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c68c6318c6318c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c68c6318c6318c626318c6e739ce739ce739ce7000"),
                (x"fffe0018c631a318c631898c6318c6e739ce739ce739ce7000"),
                (x"fffe0018c631a318c631898c6318c6e739ce739ce739ce7000"),
                (x"fffe00739c318c6318c6318c631b9ce739ce739ce739ce7000"),
                (x"fffe00739c318c6318c6318c631b9ce739ce739ce739ce7000"),
                (x"fffe00739ce70c6318c63739ce739ce739ce739ce739ce7000"),
                (x"fffe00739ce70c6318c63739ce739ce739ce739ce739ce7000"),
                (x"fffe00739ce70c6318c63739ce739ce739ce739ce739ce7000"),
                (x"ffffff8000e739ce739ce739ce739ce739ce739ce739c003ff"),
                (x"ffffff8000e739ce739ce739ce739ce739ce739ce739c003ff"),
                (x"ffffff8000e739ce739ce739ce739ce739ce739ce739c003ff"),
                (x"ffffff8000e739ce739ce739ce739ce739ce739ce739c003ff"),
                (x"ffffffffff0039ce739ce739ce739ce739ce739ce0000fffff"),
                (x"ffffffffff0039ce739ce739ce739ce739ce739ce0000fffff"),
                (x"ffffffffff0039ce739ce739ce739ce739ce739ce0000fffff"),
                (x"ffffffffffffc000001ce739ce739ce739ce000007ffffffff"),
                (x"ffffffffffffc000001ce739ce739ce739ce000007ffffffff"),
                (x"ffffffffffffffffffe000000000000000007fffffffffffff"),
                (x"ffffffffffffffffffe000000000000000007fffffffffffff"),

                -- 4_bomb_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffff8000000000000007fe94a529fffff"),
                (x"fffffffffffffffffffff8000000000000007fe94a529fffff"),
                (x"fffffffffffffff000000000000000000000000c66b5afffff"),
                (x"fffffffffffffff000000000000000000000000c66b5afffff"),
                (x"ffffffffffffc00e739ce420631b9c18c000000000000fffff"),
                (x"ffffffffffffc00e739ce420631b9c18c000000000000fffff"),
                (x"ffffffffffffc00e739ce420631b9c18c000000000000fffff"),
                (x"ffffffffff0039c39cf18c20631b9c210000001ce0000003ff"),
                (x"ffffffffff0039c39cf18c20631b9c210000001ce0000003ff"),
                (x"ffffffffff000c6210810ad6739f9cfff9ce739ce0000003ff"),
                (x"ffffffffff000c6210810ad6739f9cfff9ce739ce0000003ff"),
                (x"ffffff8000000e7210810ad6739cc6e739ce739ce739c003ff"),
                (x"ffffff8000000e7210810ad6739cc6e739ce739ce739c003ff"),
                (x"ffffff8000000e7210810ad6739cc6e739ce739ce739c003ff"),
                (x"ffffff8000000e794a5294a4739cc6e739ce739ce739c003ff"),
                (x"ffffff8000000e794a5294a4739cc6e739ce739ce739c003ff"),
                (x"ffffff8000003ff8c6318c63fffcc6e739ce739ce739c003ff"),
                (x"ffffff8000003ff8c6318c63fffcc6e739ce739ce739c003ff"),
                (x"ffffff8000000c6ffffffffe6318c6e739ce739ce739c003ff"),
                (x"ffffff8000000c6ffffffffe6318c6e739ce739ce739c003ff"),
                (x"ffffff8000000c6ffffffffe6318c6e739ce739ce739c003ff"),
                (x"ffffff80000039c318c6318dce739ce739ce739ce739c003ff"),
                (x"ffffff80000039c318c6318dce739ce739ce739ce739c003ff"),
                (x"ffffffffff00000e739ce739ce739ce739ce739ce0000003ff"),
                (x"ffffffffff00000e739ce739ce739ce739ce739ce0000003ff"),
                (x"ffffffffff00000e739ce739ce739ce739ce738000000fffff"),
                (x"ffffffffff00000e739ce739ce739ce739ce738000000fffff"),
                (x"ffffffffff00000e739ce739ce739ce739ce738000000fffff"),
                (x"ffffffffffffc00000000739ce739ce739ce000000000fffff"),
                (x"ffffffffffffc00000000739ce739ce739ce000000000fffff"),
                (x"fffffffffffffff000000000000000000000001fffffffffff"),
                (x"fffffffffffffff000000000000000000000001fffffffffff"),

                -- 5_explosion_0
                (x"ffffffb199cdada4a538c5a694a5339dad3ce739ce7bffffff"),
                (x"ffffffb199cdada4a538c5a694a5339dad3ce739ce7bffffff"),
                (x"ffffffb199ce733d6318c4eda4a53ad4e76ce739ce73ffffff"),
                (x"ffffffe739ce739b4e76b5a694a718c4e769cf39ce73ffffff"),
                (x"fffff66739ce733b5ad39e9294a529d5ad6b6739ce739cffff"),
                (x"f7bde66739cce76b5adad275a4a75ad4e73ce739ce739cb199"),
                (x"f7bde66739cce76b5adad275a4a75ad4e73ce739ce739cb199"),
                (x"739ccce739cce76b5adad27094a71a9dad9cda739e739ce66c"),
                (x"ef5999e739cce799e678c6b494a533b5ad3cdad6ce739cce6c"),
                (x"ce7399dad99ce79ce678c6a7a4a53ad4e739e6739e7339db39"),
                (x"ce7399dad99ce79ce678c6a7a4a53ad4e739e6739e7339db39"),
                (x"ce739ce733b5ad69e678c63584a5384eb56b4e73b4e79ce733"),
                (x"ce739cdad6b5ad39cf494a5294a5294eb569dad6b5ad39ce76"),
                (x"d6b539dad6b5adac4f5ad61294a5294a5389dad6b5ad6b5ad6"),
                (x"4a713b5ad6b4e7ab4d294eb49c61294a53a9dad6b5a739ced6"),
                (x"4a753b4e76b4e7ab5b494e1094a5294e3139da73b4f18c634c"),
                (x"4a753b4e76b4e7ab5b494e1094a5294e3139da73b4f18c634c"),
                (x"4a7539ce73b5ad8d5a78c25084a5294e313d6b5ab4f094a53e"),
                (x"4a756b5ad39ce78c6b5ad25094a5294e309427184eb494a53a"),
                (x"4a533b5ad34a538c2538c25384a509c2528425294eb494e138"),
                (x"c630942113c25294a5294e3094a5094e31a4a529d693ad6129"),
                (x"c630942113c25294a5294e3094a5094e31a4a529d693ad6129"),
                (x"4a529425284e309427494e128421294ce73d6a739eb139eb49"),
                (x"4a529c6b49d63094ce694e128421094253a9ce73b4e739a709"),
                (x"c613a9dad69a5294ea694a529421294a529c4f189dad39cd3a"),
                (x"4a53ab5ad69ce73d6b58c25294a709c25294ea73b5ad9ce678"),
                (x"4a53ab5ad69ce73d6b58c25294a709c25294ea73b5ad9ce678"),
                (x"d6a76b5ad6b5ad6b5a694a5294a5294a53ad4ed6b5a79cda7a"),
                (x"9ced6cce76b5ad6b5adad6b094a529d4e76b5ad6b4f339ce73"),
                (x"ce7369e733b4e76b4ed6b4d38d6b499dad6b4ed69e736b4e76"),
                (x"63339ce739ce739ce7339e138b5ad39e733b5a73ce739cce7e"),
                (x"63339ce739ce739ce7339e138b5ad39e733b5a73ce739cce7e"),
                (x"73bb9ce739ce739ce7339a71a9ce73d67399e739ce739ce72c"),
                (x"f7bb9ce739ce7339e73ad2538d6b5ac4e76b6739ce739ce739"),
                (x"ce73966739ce739b5ad6b69294a529d5ad69e739ce739ce58c"),
                (x"fffff66739ce739b5ad6b4d294a53a9dad6b6739ce739cffff"),
                (x"fffff66739ce739b5ad6b4d294a53a9dad6b6739ce739cffff"),
                (x"ffffffb199ce739b5ad6b4e78421139ce73ce739ce73ffffff"),
                (x"fffffffbd9ce739b5ad6b5ad3c613a9ce79ce739ce73ffffff"),
                (x"ffffff318cce733ccf539ceda4212842533ce739ce7339ffff"),

                -- 5_explosion_1
                (x"ce73df6739ceb494e1294a528421084253ad69299dad39e7de"),
                (x"ce73df6739ceb494e1294a528421084253ad69299dad39e7de"),
                (x"ce72cee7369a5294a7094a1084210942529c275a9ced39e599"),
                (x"9ced69ce73d2538c63094a108421084a109c6a739ced6b672c"),
                (x"b5ad6b5ad3d63094a5294a108421084a529d6b189ced39e739"),
                (x"b5ad6b4e739eb494a52842108421084a538d27189ced6b4e73"),
                (x"b5ad6b4e739eb494a52842108421084a538d27189ced6b4e73"),
                (x"b5ad6b6b5ad25294e1294a5084210842538d27189ced6b5ad3"),
                (x"9ced6b4e694a5294a7094a108421094a5294a5294ced39da73"),
                (x"4a6769dada4a5294a7094a108421384a5294a5294eb494eb53"),
                (x"4a6769dada4a5294a7094a108421384a5294a5294eb494eb53"),
                (x"4a756d6b584a538c63094a108421384a538c61294a5294a753"),
                (x"c631ac25294e3094a52842108421294a5294a7184a138c6138"),
                (x"4a5294a5294a5294a108421084210842108423184a12842709"),
                (x"4a529c6309425294a108421084210842108425294a10842708"),
                (x"4a5084a5294a1084a50842108421084210846108421094e923"),
                (x"4a5084a5294a1084a50842108421084210846108421094e923"),
                (x"4a508421084a5284a108421084210842108425294210842108"),
                (x"421084210842108421084210842108421084a5084210842108"),
                (x"42108421084210842108421084210842108421084210842108"),
                (x"421094a5284210942108421084210842108421084210842108"),
                (x"421094a5284210942108421084210842108421084210842108"),
                (x"421094a10842529c250842108421094a108421084210842109"),
                (x"423184a1084a529c250842108421084a1094a5294a10842108"),
                (x"4a5294a529421094a5084210842108425294a718c2538c2529"),
                (x"4a5294a5294a1084a5084210842108421094a1084e1294e318"),
                (x"4a5294a5294a1084a5084210842108421094a1084e1294e318"),
                (x"4a529c25294a108c2528421084210842109c25084e1294a529"),
                (x"d6b094a538c2529c63094a1084210842109461294a5294a529"),
                (x"d6b494e3094e3184a5294a1084210842109427184a5294e269"),
                (x"4a5384eb584a5294a5294a1084210842108425294a5294a678"),
                (x"4a5384eb584a5294a5294a1084210842108425294a5294a678"),
                (x"d6b534e313c25294e3094a528421084252942718c271ad4ed3"),
                (x"9ce7a4e316d2529c2538c2528421084a5284e3189cf539ce76"),
                (x"b5a739ce769a529d2538c2508421084a1084a7189dad6b5ad6"),
                (x"9cf36b5ad69e3189db094a7094210842538c6a739dad6b5a73"),
                (x"9cf36b5ad69e3189db094a7094210842538c6a739dad6b5a73"),
                (x"ce7369dad6b6b539cf494a709421094a5284e3189da79ce739"),
                (x"ce739cce769ce76d27094a52842109421084e129d5b39ce72c"),
                (x"ce739ce736b5ad84a7094a10842108421084e129d5b39ce7ae"),

                -- 5_explosion_2
                (x"fff2cce7369e3094210842108def6842109c6b18d599ef33de"),
                (x"fff2cce7369e3094210842108def6842109c6b18d599ef33de"),
                (x"fff2cce736d21084210842108bdc28421094a6739db2c6772c"),
                (x"ce58cce7339a5294a10842108bdc2842109c2673b5a79ce739"),
                (x"63199ce738d6b494a10842108bdc3b421084e3189dad9ccf39"),
                (x"9cf39ce738d6b494210842108deef7ba1084a529d4e76b5ad3"),
                (x"9cf39ce738d6b494210842108deef7ba1084a529d4e76b5ad3"),
                (x"b5a79ceb5a9eb4942108422f7bdd0842108421084ead6b4ecc"),
                (x"b5ad69eb539eb494210845c2108768425294a108c4f5ad634c"),
                (x"9ce7ad6b56d25284210845c21bdc374210842529d692842538"),
                (x"9ce7ad6b56d25284210845c21bdc374210842529d692842538"),
                (x"4a52846313c25284210845c3742377421084275a4a5294e128"),
                (x"4a50842538421084210846f68421174210846b5ac6138c6308"),
                (x"4210842109421084210842117deef742108461294a5294a529"),
                (x"4210942108421084210842021bdd1b42108425084210842108"),
                (x"421084a528421084210842361bdf77da1084a1084210842708"),
                (x"421084a528421084210842361bdf77da1084a1084210842708"),
                (x"4210842117da1084210842108086f7da1084237bba10846268"),
                (x"4210846f61da10842108423770843b421084237bdef7bda108"),
                (x"4210846f7bbdee84210845ee1084374210842108bdef7ba108"),
                (x"4210842108bdef74211bddd1708421da10842108bdc37ba108"),
                (x"4210842108bdef74211bddd1708421da10842108bdc37ba108"),
                (x"4210842108421084210846efbbdc370a1084210846efbda108"),
                (x"421084210842108421010dd1bbdee8421084210845efbda108"),
                (x"421294210842108427610a117deee842108421084210842508"),
                (x"4213a4a108421094a777bef7b4211b42108421084210842523"),
                (x"4213a4a108421094a777bef7b4211b42108421084210842523"),
                (x"4a5384a10842109d251bd86e8deee84210842108421094a51e"),
                (x"421384a529c25284a10846ef7bdc3b4210842108421094a71e"),
                (x"421094a5299eb484210846c21086f742108421294a5084231e"),
                (x"9cd284631ad25294210846c21085084210842318c6b484258c"),
                (x"9cd284631ad25294210846c21085084210842318c6b484258c"),
                (x"b5b4844e73d21094a108422fbded0842108427184eb5ad632c"),
                (x"b5b484dad6d2109d25084211b4210842109d4f5ad6b539db39"),
                (x"ce6da9dad39a5284e128422e10876842108d4e739eb539db39"),
                (x"9ced69dad69ce684a51bddc21bdd084a108c4e739e279cdb3d"),
                (x"9ced69dad69ce684a51bddc21bdd084a108c4e739e279cdb3d"),
                (x"b5ad6b5ad69ce7a4a36108421085084a5284a75a9ea79ce73e"),
                (x"ffe79b5ad6b4e7a4a2e10843b4210842538c275ab4ed9cb19e"),
                (x"fffecce739b6b49422e108437bdf6842109c275ab5b2c63bff"),

                -- 5_explosion_3
                (x"ffffef318cb25284236108421086f7da1094a75ab4f2c63bff"),
                (x"ffffef318cb25284236108421086f7da1094a75ab4f2c63bff"),
                (x"ffe79ce7399a5284211bddee1084210a10842129d6a739b273"),
                (x"b5a79cce734a52842108421010843746f68c21084eb5ad5ad9"),
                (x"b5ad9cce734a10842108422e1bdf6845ee14a529d69294ce73"),
                (x"9ced69eb494a1084211bddee1bdee845ee1ba318c61294a53a"),
                (x"9ced69eb494a1084211bddee1bdee845ee1ba318c61294a53a"),
                (x"9ced3d25294a528422e10842108437bdef7423184a52842109"),
                (x"b5a73d25294252946c2108421084210842842129c250842529"),
                (x"d6b494a52842108d8421084210842108428da129c25294a718"),
                (x"d6b494a52842108d8421084210842108428da129c25294a718"),
                (x"4a7494a5284211bbeef7b8421084210def7ba129c61294a503"),
                (x"9cf484253b42108bed17b8421084210dee10a129c21084210e"),
                (x"4a5084210842108bed17b842108421bdef70a1084a11bddf59"),
                (x"4a53bba11bddefb46c210842108437421010eef7ba101086f8"),
                (x"4a51b4211bb8421bdc210842108421421010eef70def7b86e1"),
                (x"4a51b4211bb8421bdc210842108421421010eef70def7b86e1"),
                (x"42377421170dee108421084210843746f7b0df7b0876846ee1"),
                (x"422e108421084210842108421084210842108508086fbda361"),
                (x"084370842108421084210842108421084210877b08437ba363"),
                (x"bdc37b8421084210842108421084210842108421084210deec"),
                (x"bdc37b8421084210842108421084210842108421084210deec"),
                (x"42361bdee10842108421084210842108421084210842108423"),
                (x"4211bb84210def70842108421084210842108421086e108421"),
                (x"42117bdefbbdee80842108421084210842108421bef7bddc21"),
                (x"ded08421170def708421084210842108437beef7bdd0842377"),
                (x"ded08421170def708421084210842108437beef7bdd0842377"),
                (x"4210842117ba117b84210eee10842108428422f7bed0842108"),
                (x"4210842108aa53bbdefbd8421084210defbba2f7ba10842108"),
                (x"4a5084a1084252842117b842108421ba117ba108421084213e"),
                (x"c6309425294a10842377b8437ded1708421da108421094a509"),
                (x"c6309425294a10842377b8437ded1708421da108421094a509"),
                (x"4a5294eb53c252845ef7bdef7ded1708421ba108421294e108"),
                (x"4a5294ce73c252845d17b8768421170def742529421294a67a"),
                (x"c6318d5ad34a10842117b8437bdef70dee846b184a538c4e73"),
                (x"ce593d253ad210842117b8421086f70dee8425084eb139cf39"),
                (x"ce593d253ad210842117b8421086f70dee8425084eb139cf39"),
                (x"f7bd34a5294a5294a36108421086e1bdee8421084a53ad673d"),
                (x"fffb99a5294252945c210842108421bdee842129c27539e73f"),
                (x"ffff99a10842528b842108421084210843b421294cf39ce7ff"),

                -- 6_explosion_0_0
                (x"fffffffffff3199b4d294e1294a51a9dad9b4f39ce7dffffff"),
                (x"fffffffffff3199b4d294e1294a51a9dad9b4f39ce7dffffff"),
                (x"fffffffff9ce739b4f094a5294a5389dad99cf39cb3dffffff"),
                (x"ffffffb199cce76b5a7ad4f584a53ab5ad3b4f39cb3fffffff"),
                (x"ffffffb199cce769ced6b5ad8d6b139dad3cced6cb3fffffff"),
                (x"ffffffb199ce7369eb5ad6ac94a6739dad9ce739cb19ffffff"),
                (x"ffffffb199ce7369eb5ad6ac94a6739dad9ce739cb19ffffff"),
                (x"ffffffb9cc9dad6b4e739e3484a673b5ad3ce739cb19ffffff"),
                (x"ffffffb9cc9dad3b5ad6b690842133b5ad9ce739ce7dffffff"),
                (x"ffffffb9ccb6739b5ad39a5084a7569ce799cf39cb1dffffff"),
                (x"ffffffb9ccb6739b5ad39a5084a7569ce799cf39cb1dffffff"),
                (x"ffffffffecce733b5adad2529c62769ce79b4f39f7bfffffff"),
                (x"fffffffff99dad6b5a739cd294a6769dad69e73967bfffffff"),
                (x"ffffffdad9ce736b4d38c6b09423539dad69b339cb3dffffff"),
                (x"ffffffe739ce733b69294eb5a4a5389e7339e739ce73ffffff"),
                (x"ffffffe739b5ad39cd38c271a4a529d5ad9cdad6b4e7ffffff"),
                (x"ffffffe739b5ad39cd38c271a4a529d5ad9cdad6b4e7ffffff"),
                (x"ffffffe739ce736b4e739cf494a5389dad3cdad6b673ffffff"),
                (x"fffffffbd9ce733b5a739eb094a5299dad6ccf39ce73ffffff"),
                (x"ffffffb199ce739b5ad6b61294a5294dad3ce739ce73ffffff"),
                (x"fffffffff9ce7399ce7ad6138c630944e76ce739ce73ffffff"),
                (x"fffffffff9ce7399ce7ad6138c630944e76ce739ce73ffffff"),
                (x"fffffffff9ce739ce7294a5294a7084ce79ce7396659ffffff"),
                (x"ffffffb199ce739ce6d39eb094a5294eb53ce739633fffffff"),
                (x"fffffffbccce733b4f539db094a5384eb569e739633fffffff"),
                (x"fffffffbccce736b4f539db09c63099dad39cf39ce73ffffff"),
                (x"fffffffbccce736b4f539db09c63099dad39cf39ce73ffffff"),
                (x"fffffffbd9cce76b4f539db1a9cf5ab5ad6ccf39ce59ffffff"),
                (x"ffffffb199cce76b5a739cd3a9cf56b5ad69e739cb3dffffff"),
                (x"ffffffb19d66733b5a76b6909d6a73b5ad6ce739cb1dffffff"),
                (x"ffffffffec9e7399dad39e1294a5389dad6ce73967bfffffff"),
                (x"ffffffffec9e7399dad39e1294a5389dad6ce73967bfffffff"),
                (x"fffffffff99e739cdad39eb584a509b5ad6ce739f33fffffff"),
                (x"fffffff7b99ce79cdad6b5b494a5089ce76ce7396673ffffff"),
                (x"ffffffb199cce739dad39e93a4a529d5ad69e673cb3dffffff"),
                (x"ffffffe739cce76b5ad39a753d69389dad6ce6d69e7dffffff"),
                (x"ffffffe739cce76b5ad39a753d69389dad6ce6d69e7dffffff"),
                (x"ffffffe739ce736b5ad6b6b539cd389ce73ce6d6b659ffffff"),
                (x"ffffffe739ce733b4e76b4e73c6313b5ad6ce6d6b673ffffff"),
                (x"fffff66739ce736b69339cf5a9ce739ce73ce7399e739cffff"),

                -- 6_explosion_0_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"633fffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ce739cb19dfffec67bdef33ff633d9ce736ffdce7398c633ff"),
                (x"ce739cb19dfffec67bdef33ff633d9ce736ffdce7398c633ff"),
                (x"ce739ce739cb19dce58c66739ce739ce739cb18c63339ce73f"),
                (x"ce739ce7339ce6cce739ce739ce739b67399e6d69cf39ce73e"),
                (x"ce7399ce73ce7399cf39ce739ce739b6739b6739b5b339cf2c"),
                (x"ce7399ce73ce7399cf39ce739ce739b6739b6739b5b339cf2c"),
                (x"b5a76b4e79ce733b5ad39e739ce6769ce76b4f399dad6b5b39"),
                (x"b5ad6b4e79cce76b5ad6b6733b5ad69dad6b5ad6b5a739dad6"),
                (x"d6a76b5ad6b5ad6b4e739e733b5ad39eb53b5ad6b4f539da73"),
                (x"4a676b5ad6b5ad39eb5ad5b33b5a734a5299dad6b4f56b4f09"),
                (x"9ced69ce769ce769ce739cd3ab5a73c25389ea73b4f56b6929"),
                (x"9ced69ce769ce769ce739cd3ab5a73c25389ea73b4f56b6929"),
                (x"9ce7a4eb56d631a9dad6b6938c63534eb5a9a529d6356b4d38"),
                (x"d6a7ad253ad25284e318c61294a71ac6b584a50846ad6b6929"),
                (x"d6a739eb49c2529d69294a5384a529d6b494a50842138c6129"),
                (x"9cf13d25294a53a9cf094a5384a5294a5284e1294253ad2529"),
                (x"9cf13d25294a53a9cf094a5384a5294a5284e1294253ad2529"),
                (x"9cf094a52842533d6b094a7184a5294a53a9cf5a4ce78c2528"),
                (x"9ce78c25284e313b6938c25094a5384e313b5ad69ce739eb1a"),
                (x"9ced39eb53b4e76b5a694a5284a673d4e739ce73b5a739da73"),
                (x"9ced3b5ad3b5ad6b5adad6a73b5ad6b6736b4e73b5ad6b5ad6"),
                (x"9ced3b5ad3b5ad6b5adad6a73b5ad6b6736b4e73b5ad6b5ad6"),
                (x"9ced3b5ad6b5ad6b5a76b4f369ced3cce76b6739ccf339cf39"),
                (x"ce739cce79ce7399e6739e739ce739cce739da73ce739cda76"),
                (x"ce739ce739ce739cce79ce739ce676b672ccce73ce7339ce73"),
                (x"ce6d6b4e79ce739ce739ce739ce736b6739ce739ce736b6739"),
                (x"ce6d6b4e79ce739ce739ce739ce736b6739ce739ce736b6739"),
                (x"9ced69e72cf3199ce72c63199ce736b673967b39ce739ce739"),
                (x"ce739cb19967bcc6672c63339ce7399e72cf798ccb18c63199"),
                (x"ce72cf7bd9fffeef333fffd99ce7399e73effdcef319ffffde"),
                (x"ce7fffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ce7fffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 6_explosion_1_0
                (x"ffffe667339ce769e138c4e7ad6b494a53ace739ce739cb3ff"),
                (x"ffffe667339ce769e138c4e7ad6b494a53ace739ce739cb3ff"),
                (x"ffff9cce76b5ad69a5294ea694a52842529d5a739cf39ce7ff"),
                (x"ffff9ce7399dad6d2708421084a50842538c6a73b5b39ce7ff"),
                (x"fffec66739cdad69a5284210942108425389cf5a9cf39ce7ff"),
                (x"fffffce739cdad6b4d28421294a5294a1189cf5a9cf39ce7ff"),
                (x"fffffce739cdad6b4d28421294a5294a1189cf5a9cf39ce7ff"),
                (x"fffffeb1999dad69e928421094a5284211a9eb5ace739cb3ff"),
                (x"ffffef318c9ce7a4a5294a108421084a53ad635ab672c633ff"),
                (x"fffee64e799e3094e1294a5284213ac253a9eb5ab5b3debbff"),
                (x"fffee64e799e3094e1294a5284213ac253a9eb5ab5b3debbff"),
                (x"fffff65ad69a5294e12842108421384a53ad6a739cf2c67fff"),
                (x"fffff64e76b6309c6128421084a7094a5294ea73b5ad9cffff"),
                (x"fffee66736b6b49d61294a1094a5294a5294a75ab5ad39e7ff"),
                (x"ffffdce7339eb5a9e9294a1084a5294a529c4ed6b4e739e7ff"),
                (x"ffff9cdad3d4e76b6908421084a529c6309d4f5a9cf39ce7ff"),
                (x"ffff9cdad3d4e76b6908421084a529c6309d4f5a9cf39ce7ff"),
                (x"ffffef6736b4e739e9284210842129d63094a5299dad9cf7ff"),
                (x"ffffef6739b5ad39eb58c2508421084a5294a718b5a79cb3ff"),
                (x"ffffd66733cdad3d6b094a508421094a5294a7189e739cb3ff"),
                (x"fffee66733b5ad6b4f094a108421084e3094eb189db39ce7ff"),
                (x"fffee66733b5ad6b4f094a108421084e3094eb189db39ce7ff"),
                (x"ffffdce739cce739db494a508421084a5294ce739dad9ce7ff"),
                (x"fffecce739cce7a9cf494a509421094a5294ced6b4ed9ce7ff"),
                (x"ffff9cb1999dad3d6938c250842108425294ea739ced39e7ff"),
                (x"fffff63193b5ad3d2538c2108421084253ad6b18d5ad39e7ff"),
                (x"fffff63193b5ad3d2538c2108421084253ad6b18d5ad39e7ff"),
                (x"fffffee7369ce734a7094a508421184e31ad4f18d5ad39e7ff"),
                (x"ffffef31999e3094e1294e928421184a53a9ea73ce739ce7ff"),
                (x"fffec67bccb6b494a5294a528421094a5294ead6ce739ce7ff"),
                (x"fffff731999eb53d25084210842109c25294ead6b6739cffff"),
                (x"fffff731999eb53d25084210842109c25294ead6b6739cffff"),
                (x"fffff731999a533b69294a1094a509c25339ced69e72c67fff"),
                (x"ffff373193b253ab4d294a1094a5384e3169ead6b658e77bff"),
                (x"fffec667369a533b4f494a108421094e31ac6273b5b2c633ff"),
                (x"ffffdcdad39dad69e3484210842108425384ea73cced9ce7ff"),
                (x"ffffdcdad39dad69e3484210842108425384ea73cced9ce7ff"),
                (x"ffff99dad6b4e73d25294a10842108425294e273ce739ce7ff"),
                (x"ffff99e7399ce7a4a5094a108421084a5384ead6b5a79cb3ff"),
                (x"f7999ce733c63094a10842108421094e3094ced6b5ad39b3ff"),

                -- 6_explosion_1_1
                (x"f7bfffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"f7bfffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"633fffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ce739eb193fffecf7ff9cb3aeef7decf7aeffdcef7fec6673e"),
                (x"ce673cb18e739ccf7599ce72c633dece72c6318cf772c6672c"),
                (x"ce736b672c6319e6658c66739ce739b67399da7363339ce679"),
                (x"ce736b672c6319e6658c66739ce739b67399da7363339ce679"),
                (x"9cf369dad3ce72ccda79ce7339cf369ce76b5b3966739ce6d3"),
                (x"c62769ce769ce769ced39e736ce6d6d4e76b4e739cf39cced3"),
                (x"c6273b25294eb5ac4ed6b4e76b5ad39eb5ac27189dad6b5ad3"),
                (x"c6273b25294eb5ac4ed6b4e76b5ad39eb5ac27189dad6b5ad3"),
                (x"4a753b4e7a9ce694ce739ea769ce73b6b494a529d5ad6b5ad6"),
                (x"4a53a9dad6b6b494a75ad4e76d6a73b4e7ac25294ced39ea73"),
                (x"42129c4e73d2529c253ad4ed3d6b5ad6b58c63184ea694a538"),
                (x"42109d6b494a1094e1294eb58c6349425294a5294a5294e129"),
                (x"42129425294a1094a718c25294a70842529421294a10842138"),
                (x"42129425294a1094a718c25294a70842529421294a10842138"),
                (x"421084210842109d25094a5284a52842108421294210842353"),
                (x"4210842108421094a108421084210842108421294212842273"),
                (x"42108421094a1084210842508421084210942108425294a13a"),
                (x"42108421094a1084210842108421084a5294a108425284253a"),
                (x"42108421094a1084210842108421084a5294a108425284253a"),
                (x"4210842109421084210842108421094a529c2529425284213a"),
                (x"4a508425384a529c6108425084a5094a5294e35a4212842109"),
                (x"4a52842529c63094a508425294a53ac25294a7184a12842109"),
                (x"c61294e3184a5294e1294a5384a538c25294a5294a1094a529"),
                (x"c61294e3184a5294e1294a5384a538c25294a5294a1094a529"),
                (x"4a709c6b569a529d6b494a5294a5294a5294eb5ad6b18c613a"),
                (x"4a5294e3139a5299eb494a5294a529d63094ea73d4e739e359"),
                (x"9cf58d631a9eb5ad4f5ad4e7a4a5299ce69d6b5ac6a739ead9"),
                (x"b5ad39ce76b5ad69e3139da78c6309d5ada9cf5ad6b5ad4e79"),
                (x"b5ad39ce76b5ad69e3139da78c6309d5ada9cf5ad6b5ad4e79"),
                (x"b5ad9cdad69dad9ceb539da739ced39dad6b4ed6b66739da79"),
                (x"b5ad99dad9ce739cdad39ced6ce6d69ce76b4ed6ce6739da79"),
                (x"b5a79b672cce739cdad6b5ad9ce676cce76b6739ce739ce739"),
                (x"9cf39cb18e66739cce739e739ce739cce73cb3bd66739ce739"),
                (x"9cf39cb18e66739cce739e739ce739cce73cb3bd66739ce739"),
                (x"63199cb19effff9ce739ce7396319dce739ffdce63339ce72c"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 6_explosion_2_0
                (x"ffd8ccce769e3094250846f77ded084a53a4a75a9dad6b67df"),
                (x"ffd8ccce769e3094250846f77ded084a53a4a75a9dad6b67df"),
                (x"ffd99cce769eb53c250842361bdd084a53a4a75ad4ed6b4d9f"),
                (x"fff39cce76b4e73d250842117bdc37421084275a9cf56b673f"),
                (x"ffd8ccdad6b6b49c210842377bdee1ba108421084e356b659f"),
                (x"fffdd65ad69e3094a1084211bbdc3b42108421084a676b31df"),
                (x"fffdd65ad69e3094a1084211bbdc3b42108421084a676b31df"),
                (x"ffffff4e76b6b494a10842117bdc28421084275a9dad6b31df"),
                (x"ffffff6733b5ada4210842108dec284210842129d5ad9cb3ff"),
                (x"ffd9eee736b5ad3421294a108422fbda10846b5ad5ad9cfbff"),
                (x"ffd9eee736b5ad3421294a108422fbda10846b5ad5ad9cfbff"),
                (x"ffd2cce736b4e73c2128422fb4211bba108c4ed69dacc67b3f"),
                (x"ffd13cdad69e309421284202108421bef684275a9ea6c6667f"),
                (x"ffd19cce739a5294210842021084210dee842129d4e79ce73f"),
                (x"ffd036319a9ce7a4e108422f7bdc37bef684a1089da6c6659f"),
                (x"ffd1ad6733d5ad3d612846c370843b421084a673b4f39ce7df"),
                (x"ffd1ad6733d5ad3d612846c370843b421084a673b4f39ce7df"),
                (x"fff19b6733b5ad34a528422e1bdee842109426d6b5ad9ce7df"),
                (x"fff19ce7399dad3c2108422f7def684252944ed69dad9cb1df"),
                (x"ffd19ce739cdad6d21294a117ded0842538d4ed69dad9ce59f"),
                (x"fff19ce739cce7a4212842108bdee8425294ce73d4e79ce73f"),
                (x"fff19ce739cce7a4212842108bdee8425294ce73d4e79ce73f"),
                (x"fff59b5ad39eb48425294a361bdef7da1094235a4ea79ce73f"),
                (x"fff0ccdad3b5ac94a10842108bdc21bef684a1299ce79ce73f"),
                (x"ffd3dce733b4e7a4210842377bdf77da1084235ab5b39ce73f"),
                (x"ffdddce733b6b494210842361bdd084210842673b4e79ce73f"),
                (x"ffdddce733b6b494210842361bdd084210842673b4e79ce73f"),
                (x"fffff66736b4e69421084237b42108421084235a9e72c65b3f"),
                (x"ffffff7bd9b5ada42108421084211bda1084a673d633decfff"),
                (x"fffcc63193b4e734a5294a108bdc3742108c4e73d266c63bff"),
                (x"fffccf6733b6b494a5284211bbdefb42108d4f5ab4f539b3bf"),
                (x"fffccf6733b6b494a5284211bbdefb42108d4f5ab4f539b3bf"),
                (x"fff39cce769a5384210842108bdef742108c5a739cf539e59f"),
                (x"ffe799dad69ce734a12842108bdc3b421084ce739ce76b599f"),
                (x"ffe76b5ad69dad34a5094a108bdc28425294a5299dad6b5b3f"),
                (x"fff339dad3d5ada4a5084211b086fb4e3094a5299e679ccf3f"),
                (x"fff339dad3d5ada4a5084211b086fb4e3094a5299e679ccf3f"),
                (x"fffd9ce7334ce739e92842101bdefb425294a508d6739ce73f"),
                (x"fffd9ce7339eb53b4f494a2e1bdf6842538421084da79ce73f"),
                (x"ffe76b4e76b4e73b4f08422e84210842538c25084a539ce73d"),

                -- 6_explosion_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"9cfdecce73cfbdeffdc94e35842318421084258cfffcc6658c"),
                (x"b5b399dad9cb18cfffbdeb339ce739d0c799b3defffac6672c"),
                (x"b5b399dad3cfbccf3339ce6d9ce736d3199ce7bdf7999ce739"),
                (x"9cf39b5ad69e72cf6739cdad9ce739cb193b6739cced6b4e73"),
                (x"9cf39b5ad69e72cf6739cdad9ce739cb193b6739cced6b4e73"),
                (x"b5a739dad6b4e73cda739ce79ce7339eb53b5ad69dad6b5ad6"),
                (x"b5a69d4e739dad6b5ad6b5a79ce676d4e739dad6b5a76b5a73"),
                (x"9cf53b5ad34eb53b4f539db53b5ad6b4e69c4ed6b6b1ad4f58"),
                (x"9cf53b5ad34eb53b4f539db53b5ad6b4e69c4ed6b6b1ad4f58"),
                (x"9ce73d4e73c2533d253ad251ab5a739eb494ce73d25294ce69"),
                (x"b5ad34a529425294210842508d6b09d25284610842538c6b08"),
                (x"9ce7a4a52842529421084212842109c6308421084210842529"),
                (x"c6349421094252942108421294a5094a1084a5294210842108"),
                (x"42128425284210942108421284a50842108421294210842108"),
                (x"42128425284210942108421284a50842108421294210842108"),
                (x"421084210842108421084210842108da10842108421084211b"),
                (x"bdee8421084210846f7bda368422f70dee10dd084211bda37b"),
                (x"42021da10846f6846c37ba028bdee1bdee10ed0845f77bdc37"),
                (x"422f70def7bdef7422f7bdef7def770dee10a108ddef7bdefb"),
                (x"422f70def7bdef7422f7bdef7def770dee10a108ddef7bdefb"),
                (x"42377b8421bdee14211bd86f742377084210a2f708437b8508"),
                (x"4211bda11bbef77da117b86e842108ddee10ef7b423610dd08"),
                (x"421084a10842108da11bddf684210845ee1bdf7b42117ba129"),
                (x"4a529c2528421084210846d094a52846f77da1084210842129"),
                (x"4a529c2528421084210846d094a52846f77da1084210842129"),
                (x"c63094a528421084210842129c61294210842108421084235a"),
                (x"c61094a529c6b584a10842509d69084a528461084210842129"),
                (x"4a5094a533b4e734a128421139ce694a1084cf5a4250842529"),
                (x"421084a5339eb539ea7ad2753b5ad69a109d5b5a4e90846b5a"),
                (x"421084a5339eb539ea7ad2753b5ad69a109d5b5a4e90846b5a"),
                (x"4a53a9ce739dadad4ed6b4d3a9ce76b4e7a9cf5ad4d294cf53"),
                (x"4a6d9cdad39ce69c6676b4f53b5ad69dad3d5ad6b5938c4e76"),
                (x"4a6799dad3d6b53ce679cce73b5ad6cce739dad6b5a7ad6ad6"),
                (x"ce739cdad69ce6ceb339ce739ce739cb19963339cdad6b5ad6"),
                (x"ce739cdad69ce6ceb339ce739ce739cb19963339cdad6b5ad6"),
                (x"ce7399dad6cb18e9db39ce739ce599ce739cfbde63199ce679"),
                (x"ce739ce72c677bffe739ce739631def31999e7fffb9cc6659e"),
                (x"f7bfffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 6_explosion_3_0
                (x"b5a73b5ad6b5ad69a508421084210842529d2108426739e58c"),
                (x"b5a73b5ad6b5ad69a508421084210842529d2108426739e58c"),
                (x"633399ce769ce73d251bddc3b4211bda10842108421294cf39"),
                (x"ef7cc9dad34a108423610843b422e1ba108425084a53ad673f"),
                (x"fffecce7334a108422b7b86f7bdc21bef694a508c6b539e7ff"),
                (x"ffffdce73a4a5284210845f61084210dee842508c4ed39e7ff"),
                (x"ffffdce73a4a5284210845f61084210dee842508c4ed39e7ff"),
                (x"ffff9b673a425294a50845c21086e10843b42529c5b39ce59f"),
                (x"fffecb5ad3425284a53bddc3bbdee10843742129c4ed39e7ce"),
                (x"ffff3b5ad34e3094a108406fb08421bdee8421294ced6b658c"),
                (x"ffff3b5ad34e3094a108406fb08421bdee8421294ced6b658c"),
                (x"ffff6b5ad34a5384a10846c21bdc21ba10842108d5ad6b5a79"),
                (x"632d3d4e7ac25294a11bddc21bdf61ba11b421084ce739e739"),
                (x"ce673d25294a10842117b8421ded17084374210842759ce73f"),
                (x"ce7369a5294210842117b842108421ba108421084ead6b5bff"),
                (x"d6b36d2538421094236108421bdc370ef68421294ead6b5bff"),
                (x"d6b36d2538421094236108421bdc370ef68421294ead6b5bff"),
                (x"ce7369eb53c25294236108421bdc28def6842129c4ed6b5bff"),
                (x"b5b39b5ad6d21094211bd86f7bdef742108425294eb539dbff"),
                (x"63279b5ad3c25294eefbddd0842377da108425294eb539cf3d"),
                (x"ce6769dad6d21084236842108deefb421084210846a76b658c"),
                (x"ce6769dad6d21084236842108deefb421084210846a76b658c"),
                (x"ce739cce76d210842108422fbbdef742528421084ce79cb199"),
                (x"d6999cdad3d25284211bddc210876142529421084ce739f99f"),
                (x"ffff9cdad64a1084236108421def61da1084a52946a739cfff"),
                (x"ffff99ce73421084210845efbdeee1ba10842718d62739e7ff"),
                (x"ffff99ce73421084210845efbdeee1ba10842718d62739e7ff"),
                (x"ffffac2528425284210846f7708421ba1094e1294e2739e59f"),
                (x"fffe94a52842108422f7bdee108437da1094e3184cf39ce739"),
                (x"ffff39ce7a4210842361086e1bdefbda10842529d4ed39e739"),
                (x"ffff6b5ad3c25284236108421ded17ba108421084dad39e72c"),
                (x"ffff6b5ad3c25284236108421ded17ba108421084dad39e72c"),
                (x"18d96b5ad69a528422e1084210843b0ef684210844ed6b33de"),
                (x"d6bb6b4e76d252842117b84210843b0ef68421084da76b7bcc"),
                (x"ce7369ce73c2108ddee10842108437ba1084210844e739b3ff"),
                (x"ce733b5ad84a108d84210eee1084210dee84210846279cf7ff"),
                (x"ce733b5ad84a108d84210eee1084210dee84210846279cf7ff"),
                (x"f7bb9b4e694252846c210dc3b084210def7421294ce6c63bff"),
                (x"ffdcccce69d2528422e10defb420374210842129c6a79ce7ff"),
                (x"fffeceb19a9a528422fbda37b422f74210842129c27139dbff"),

                -- 6_explosion_3_1
                (x"ffffece73a1ffffffffffeb39632d9d673967ffffffffff596"),
                (x"ffffece73a1ffffffffffeb39632d9d673967ffffffffff596"),
                (x"ffdddce73d67fffffffffb3339cf39ce733b7ffffffffffb33"),
                (x"631999dad6b5ad34eb39ce736ce736b5ad39da73667ac63333"),
                (x"ef736b4e76b5ad34e279ce733b5ad3d4e7ad5ad6b5b39cce76"),
                (x"63273b4e73b5ad34a676b5a76b5ada4a5299dad6b6739cda76"),
                (x"63273b4e73b5ad34a676b5a76b5ada4a5299dad6b6739cda76"),
                (x"d6929c4e76b4e7a42276b4ed69ced3c2529d4e739eb539ced6"),
                (x"9cf484e31a9e308421094eb5ac635842109c2529421294a676"),
                (x"4a529421094a52842508425084a509421084a7184a52842276"),
                (x"4a529421094a52842508425084a509421084a7184a52842276"),
                (x"42108421084210842108421084a5294a1084e1294250842276"),
                (x"42108def684210842108421084a508421084a5294a50842353"),
                (x"4211b0dee8421084210842108ded0842108421084a50842129"),
                (x"bdee10dee8bef7bba11bda11bbdd1bda108421084a115aed08"),
                (x"dec210843708421ba1010ed08def610def7da108da117b8768"),
                (x"dec210843708421ba1010ed08def610def7da108da117b8768"),
                (x"422f7d842108421beee10dd08bdc2108421bec21bdee1086e8"),
                (x"deee1b842108437beee1086e8422e108421086f708777b8428"),
                (x"def7b08421084210df6108768422e1084210877bd8437bef68"),
                (x"42101084210ef770877bd86fb422f7b843bbdc21b8437ba108"),
                (x"42101084210ef770877bd86fb422f7b843bbdc21b8437ba108"),
                (x"bdc21084210a117086fbdeef7deee108428d8421bdc210dd08"),
                (x"bdee10defbddefbb8421086fbbdee8b8437084210842108768"),
                (x"421010dee10defbddefbda108ded1b0dee1bdef708437bdf68"),
                (x"42117ba11bda10842108425284211bda101422f7086fbda109"),
                (x"42117ba11bda10842108425284211bda101422f7086fbda109"),
                (x"4211742108421084a508425084210842117da108bed094a109"),
                (x"4210842108421084a5094a108421084210842108421094a11a"),
                (x"421084210842109c61294a1084a5284210842108425294a508"),
                (x"4a5294210842109c27094a1084a5294a108421294a50842108"),
                (x"4a5294210842109c27094a1084a5294a108421294a50842108"),
                (x"c6309421094253a4a748425284a5384a5284e929c6318c2508"),
                (x"4a753c4e769dad39e31ad4e7ad6b53d6b499da739da7ad2509"),
                (x"c62739ce73b5ad6cce739ce73d6b56b5ada9dad6b66dad2533"),
                (x"9cf2ccce76b4e73cce739cf369ce76b5ad99dad69e6739e933"),
                (x"9cf2ccce76b4e73cce739cf369ce76b5ad99dad69e6739e933"),
                (x"b5b2eeb19e66739ce7339f9999ced6b5ad9cdb39ce739ce679"),
                (x"fffffffffef6739cb3fffb18cce7ffffff9ccd8cf33fffe72c"),
                (x"ffffffffecf3199cfffffff2cef7fffffffce58c77ffffff2c"),

                -- 7_explosion_0_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffef332cce739cfffffffffffffffffff"),
                (x"ffffffffffffffffff39ce739ce739ce73ffffffffffffffff"),
                (x"ffffffffffffff9ce739ce739ce739ce739cb3ffffffffffff"),
                (x"ffffffffffffff9ce739ce739ce739ce739cb3ffffffffffff"),
                (x"fffffffffffe739ccf39ce739ce7339e739cb18cffffffffff"),
                (x"fffffffffff6739cdb39ce739ce7339dad3ce739cfffffffff"),
                (x"ffffffffff667399e739ce739ce6d6b5ad3ce739cfffffffff"),
                (x"ffffffffff667399e739ce739ce6d6b5ad3ce739cfffffffff"),
                (x"ffffffffffce7339e679ce679ce6d39ce79ce739cfffffffff"),
                (x"ffffffffecce739cdb39ce6739cf33cce73ce739cb3fffffff"),
                (x"ffffffb18cce739cce79ce6d6b5ad6cce73b5b39cb1dffffff"),
                (x"ffffffe739ce739cce76b66d6b5ad6b5ad6b4f39ce7bffffff"),
                (x"ffffffb199ce739ce676b4f53b5a73b5ad6b4f39ce59ffffff"),
                (x"ffffffb199ce739ce676b4f53b5a73b5ad6b4f39ce59ffffff"),
                (x"ffffffe739ce733ccf56b6929c6133b5ad69e739ce59ffffff"),
                (x"ffffffe739ce7399da76b69384a53a9dad3ce739ce7fffffff"),
                (x"ffffffe739ce739cced39e1294a7494eb53ce739ce7fffffff"),
                (x"fffffffff9ce739ce6d39e1294a753d6b539cf39ce7bffffff"),
                (x"fffffffff9ce739ce6d39e1294a753d6b539cf39ce7bffffff"),
                (x"fffffffff9cdad3cdad39a53a9ced6b5ad39dad6b67bffffff"),
                (x"ffffffe7399dad6cdadad253a9cf53b4e7a9da739e59ffffff"),
                (x"ffffffe7399dad6b5ad39e933d6b1a9ce769e739ce59ffffff"),
                (x"ffffffe739cdad6b5adad6b53d6a7a4ce76ce739ce59ffffff"),
                (x"ffffffe739cdad6b5adad6b53d6a7a4ce76ce739ce59ffffff"),
                (x"ffffffb199ce736b5ad39e273d6a739dad69e739ce73ffffff"),
                (x"fffffffffece739b5ad6b4e784a5339ce76b6739ce7fffffff"),
                (x"ffffffffeef3199cced6b5b094a7139ce76b6739cb3fffffff"),
                (x"fffffffbdef7bd9cced6b4d294a713d4e739da73cf7dffffff"),
                (x"fffffffbdef7bd9cced6b4d294a713d4e739da73cf7dffffff"),
                (x"fffffffbdece7399ced39e129d6b5a9ce739dad6cfbdffffff"),
                (x"fffffffbccce733b4ed6b6938d6b18d4e739cf39cb19ffffff"),
                (x"ffffffb9ccce733b5a739cf58d6b5ad6b5a9ce73ce73ffffff"),
                (x"ffffffb9cc66733b4f539db49d6b58c6b5a9ce7367bbffffff"),
                (x"ffffffb9cc66733b4f539db49d6b58c6b5a9ce7367bbffffff"),
                (x"ffffff7bdece739b5a76b4f094a753d6b58d4e73cb19ffffff"),
                (x"ffffffb9ccce7339ce76b4f49c635ad4e7ad4e73ce73ffffff"),
                (x"ffffffb9ccce73964e739cf5ac635a9ce739cf39f7bbffffff"),

                -- 7_explosion_0_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffefffffffffffffffffffffffffffffffffffffffffffff"),
                (x"739de739def7bdffb339ce7ffce7396672cfffffffffffffff"),
                (x"739de739def7bdffb339ce7ffce7396672cfffffffffffffff"),
                (x"6319e6318cf7bcef6739ce739ce739ce72c67fffffffffffff"),
                (x"ce73966739cfbdece7339cf39ce739ce739ce58cf7ffffffff"),
                (x"ce739ce739cfbccce6d6b5ad9ce739ce739ce739ce7fffffff"),
                (x"ce739ce739cfbccce6d6b5ad9ce739ce739ce739ce7fffffff"),
                (x"ce6799ce73ce739cdad6b5a79ce733ce739ccf39ce73ffffff"),
                (x"63276b5ad69e739b5ad6b6739ce679ce739cce73ce73ffffff"),
                (x"9ce769dad39ce73b5ad6b5ad99ced3cce73b6739b4f3ffffff"),
                (x"9ce73d4e76b5ad6b5ad6b5ad6b5a7a9ce73ccf39ce739cffff"),
                (x"9ced69ce769dad6b4f539ea739ced6b5ad9ce739ce739cfbff"),
                (x"9ced69ce769dad6b4f539ea739ced6b5ad9ce739ce739cfbff"),
                (x"9ce73b4e7ac4e769e35ad2538c635a9e739ce739ce739cb3ff"),
                (x"d6b58d6b494a5389cf494a5294a529d5ad69cf39ce739ce7ff"),
                (x"d69294e3184a529c4e739eb494a7099dad69e739ce739cb3ff"),
                (x"c6309d6b5ad25294eb5ad4e694a538b5ad69e739ce739ce7ff"),
                (x"c6309d6b5ad25294eb5ad4e694a538b5ad69e739ce739ce7ff"),
                (x"d6b5ad6b58d63184ce78c6adad69299dad6cdad6ce739ce7ff"),
                (x"d6b53c6b58d4e739cf5ad4ed34a7539dad69ced69cf39ce7ff"),
                (x"9cf5ac6b5a9eb539cd339dada4a676b5ad9cced69cf39ce7ff"),
                (x"9ce7ad6b539ce739da739cedad6ad6b5ad39ced6b6739cffff"),
                (x"9ce7ad6b539ce739da739cedad6ad6b5ad39ced6b6739cffff"),
                (x"9cf58d6b539ce76b5ad6b6a739ce76b5ad39e6739e73ffffff"),
                (x"9cf5a9ce739ce76b4f339ce73ce733b5ad6ce739ce73ffffff"),
                (x"9ce739ce73b5ad9ce739cdad3ce7399ce76ce739cb19ffffff"),
                (x"ce6739ce79b4e79ce739cced9ce739ce739ce739cb3fffffff"),
                (x"ce6739ce79b4e79ce739cced9ce739ce739ce739cb3fffffff"),
                (x"f7b3966739ce739ce739cced9ce739ce739ce739cfffffffff"),
                (x"f7b2cf672cf77acce739ce739ce739ce72c67fffffffffffff"),
                (x"ef72cee72cf7bdffe58c633bdfffec677aefffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_0_2
                (x"fffffff7bef67339ce739eb58d6b539ce7366739cb1dffffff"),
                (x"fffffff7bef67339ce739eb58d6b539ce7366739cb1dffffff"),
                (x"ffffffe739cce73d6a7ad6b584a753b4e739cf39cb1dffffff"),
                (x"ffffffb18ccce73d635ad4f494a713b4e76b6739cfbdef7fff"),
                (x"fffffff7be64e739eb58c635a4a7569eb53b4f39631dffffff"),
                (x"ffffffe739cce739eb5ad6b5ac63539ce76b4f39cb1dffffff"),
                (x"ffffffe739cce739eb5ad6b5ac63539ce76b4f39cb1dffffff"),
                (x"ffffffb18cce7339ce7ad631ac613ab5ad3b4f39cb3dffffff"),
                (x"fffffffbdecdad69ce739eb5a4a5389dad39e739cfbdffffff"),
                (x"fffffffbddcce769ce7ad4f094a533b5ad3ce7def7bdffffff"),
                (x"fffffffbddcce769ce7ad4f094a533b5ad3ce7def7bdffffff"),
                (x"ffffffffecce739b5a739cf094a716b5ad3ce58cf3bfffffff"),
                (x"fffffffff9ce739b5a739cd29c6273b5ad6b6739cfbfffffff"),
                (x"ffffffe739ce7399dad39ce7a9ce789dad6b5b39ce59ffffff"),
                (x"ffffffb199ce739cda694ea7a9cf5ad5ad6b5ad6ce73ffffff"),
                (x"ffffffb199ce7399da739eb1a9cd3a9dad6b5ad69e73ffffff"),
                (x"ffffffb199ce7399da739eb1a9cd3a9dad6b5ad69e73ffffff"),
                (x"ffffffb1999ce769ea76b4f53d6929d5ad6cdad69e73ffffff"),
                (x"fffffff7b9b5ad69ced6b5ad3d69299dad6cced6ce7fffffff"),
                (x"fffffff7b9ce7339cf5ad4f494a5389dad9ce739ce7fffffff"),
                (x"fffffffff9ce739ccf494a7494a5389dad3ce739ce73ffffff"),
                (x"fffffffff9ce739ccf494a7494a5389dad3ce739ce73ffffff"),
                (x"fffffffff9ce739cced39e929c613ab4e769e739ce73ffffff"),
                (x"ffffffb199ce7399dad6b4d384a53ab6b53ccf39ce73ffffff"),
                (x"ffffffb199ce733b5ad6b4e769cf53b4e79ce739ce59ffffff"),
                (x"fffffff7b9ce733b5ad6b5ad6b5ad9b4e73ce739ce73ffffff"),
                (x"fffffff7b9ce733b5ad6b5ad6b5ad9b4e73ce739ce73ffffff"),
                (x"ffffffb9ccce736b4e79cdad6b5ad9cce73ce739cb19ffffff"),
                (x"ffffffffecce739cce79ccf339ce79ce736ce739cb3fffffff"),
                (x"ffffffffffce739ce6739ced9ce679cce799cf39cfffffffff"),
                (x"ffffffffffce739cced6b5ad9ce739ce7399e73967ffffffff"),
                (x"ffffffffffce739cced6b5ad9ce739ce7399e73967ffffffff"),
                (x"ffffffffffce739cced39cf39ce739ce736ce739f7ffffffff"),
                (x"fffffffffffb18cce7339cf39ce739ce733ce739ffffffffff"),
                (x"fffffffffffffecce739ce739ce739ce739ce7ffffffffffff"),
                (x"ffffffffffffffffff39ce739ce739ce73ffffffffffffffff"),
                (x"ffffffffffffffffff39ce739ce739ce73ffffffffffffffff"),
                (x"fffffffffffffffffff9ce7396332cf7ffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_0_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffbbac633ffef7ac63199fffdef333deb33d"),
                (x"ffffffffffffffffbbac633ffef7ac63199fffdef333deb33d"),
                (x"fffffffffffffff63339ce739ce739ce739cb3bdf333ef333e"),
                (x"ffffffffffce739ce739ce739ce6d3ce739ce739ce72c6673e"),
                (x"ffffffffecce739ce739ce739ce6d3ce739ce673b66739ce79"),
                (x"ffffffffecce739ce739ce739ce6d3ce739ce673b66739ce79"),
                (x"ffffffb18cce739cda739e7399ced6ce739ce6d6b4e739ce73"),
                (x"ffffffe739ce739cdad6b4f399ce739e733b5a739ce739eb53"),
                (x"ffffffe7399ce799ced6b5a739ce7ab5ad6b5a739cf5ad6353"),
                (x"fffffce739b5ad39ced6b5adad6ad39ce769ce739cf5ad6a73"),
                (x"ffff9ce7339dad3ce6d6b5a69d6ad69a5339cf5a9eb58c6b53"),
                (x"ffff9ce7339dad3ce6d6b5a69d6ad69a5339cf5a9eb58c6b53"),
                (x"ffff9ce7339dad39dad39cf499ced3d6b539ce73d6358c4f5a"),
                (x"ffff9ce739cdad6cdad39a53ad6adac4e734e318d635ad6b5a"),
                (x"ffff9ce739ce7399dad6b61294a673d6b5a4a529d6b5ad2718"),
                (x"fffecce739ce7399dad39a7094a75a9ce73c25294e3094a53a"),
                (x"fffecce739ce7399dad39a7094a75a9ce73c25294e3094a53a"),
                (x"ffff9ce739ce7339dadad25294a5294eb539e1294a75ad635a"),
                (x"fffecce739ce739ce7339eb58c6129d6b589da73c6a76b4e73"),
                (x"ffffece739ce739ce6d6b5ad39ce7a9eb53b5ad69da739dad3"),
                (x"fffffce739ce733cce739ea76b5ad6b5ad6b5ad6b5a7ad4e73"),
                (x"fffffce739ce733cce739ea76b5ad6b5ad6b5ad6b5a7ad4e73"),
                (x"ffffffe733b6739b4e79cced3ce6d6b5ad6b4e739ced39da73"),
                (x"ffffffe739cce73ce739ce679ce739b5ad6b67399dad6b5a6c"),
                (x"ffffffe739ce733ce739ccf39ce676b5ad6ce739cce739e679"),
                (x"fffffffff9ce739ce739ce739ce6d6b5ad9cb3dece739ce739"),
                (x"fffffffff9ce739ce739ce739ce6d6b5ad9cb3dece739ce739"),
                (x"fffffffffff3199ce739ce739ce7339e739cfbdece72c66739"),
                (x"fffffffffffffff63339ce739ce739ce739f3bdef318c6798c"),
                (x"ffffffffffffffffb32c66739ffff9ce72cfffdef79ce779ce"),
                (x"fffffffffffffffffffffffffffffffffffffffffffffffbff"),
                (x"fffffffffffffffffffffffffffffffffffffffffffffffbff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_1_0
                (x"ffffffffffffffffffffffffffff5a9eb539cf39ffffffffff"),
                (x"ffffffffffffffffffffffffffff5a9eb539cf39ffffffffff"),
                (x"fffffffffffffffffff9cce796319ecfffffffffffffffffff"),
                (x"ffffffffffffffffff39cdad3ce739ce73ffffffffffffffff"),
                (x"ffffffffffffbdece6739dad6b5b39ce73963bffffffffffff"),
                (x"fffffffffffb19ece6d6b5ad6b5a73ce739cb3bdffffffffff"),
                (x"fffffffffffb19ece6d6b5ad6b5a73ce739cb3bdffffffffff"),
                (x"ffffffffffeb199ce6739ced39ced6b6739ce58cf7ffffffff"),
                (x"fffffffff9cb199ce6739dad69ced6b5ad9ce739ccffffffff"),
                (x"ffffffb193b6739ccedad4ed6b5ad6b5ad99dad6b4d9ffffff"),
                (x"ffffffb193b6739ccedad4ed6b5ad6b5ad99dad6b4d9ffffff"),
                (x"ffffffe739b4e76b4e7ad6ad69ce739ce739dad6b4f3deffff"),
                (x"ffffffe7399dad6b6b58c6a739cd3ac25389dad69e72c67bff"),
                (x"fffffce7339dad69a53ad6b53d69294eb5ad4ed6b4f39cb3ff"),
                (x"fffeccdad3cce76d2538c4e7a4a529d5ad3c6ad6b4f39cffff"),
                (x"ffff9cdad3ce7369eb494eb094a53ad5ad3c6ad6b4ed6b7fff"),
                (x"ffff9cdad3ce7369eb494eb094a53ad5ad3c6ad6b4ed6b7fff"),
                (x"ffff9ce7339ce7ad6b094a5284a538c6b494ead6b5ad39e7ff"),
                (x"ffff9ce733b4e694e938c25284a7094a53ac4ed6b5ad9ce7ff"),
                (x"ffff9cce769ce784a5294e128421294e313b5ad6b5a79ce7ff"),
                (x"ffff9cdad6b4e784a538c252842109c253ab4ed6b4f39ce7ff"),
                (x"ffff9cdad6b4e784a538c252842109c253ab4ed6b4f39ce7ff"),
                (x"ffff9ce736b5ada4a5294a10842109c2529d635ab5b39ce7ff"),
                (x"ffff9cce73d6b53d4f494a10842109c2538d69299db2c633ff"),
                (x"ffff9cdada9dad6b5b494a70842109c2533b4f5ad5b3deffff"),
                (x"ffff9cce7ad4e73d61294a52842109c253a9ced69da79cffff"),
                (x"ffff9cce7ad4e73d61294a52842109c253a9ced69da79cffff"),
                (x"ffff9cce78c4e7a4a538c2508421294a529c6ad6b5a79cb3ff"),
                (x"ffff9cce739ce694a538c25284212846309d4ed6b4f39ce7ff"),
                (x"fffffce733b4e694a5294a5284210842538d4f39ce739cffff"),
                (x"fffff667399dad3d25294a108421084e3189ce73cb199cffff"),
                (x"fffff667399dad3d25294a108421084e3189ce73cb199cffff"),
                (x"fffecce733b5ad6b6938c2508421094a5389ead69e599ce7ff"),
                (x"ffff9ce733b5ad69e9294a108421094a53ab4f5a9e72c633ff"),
                (x"ffff9cce76b5ad69e1294a108421094a533b4d29d659ef33ff"),
                (x"ffff9ce736b5ad6b692842108421094a533b5a739cd9ef77ff"),
                (x"ffff9ce736b5ad6b692842108421094a533b5a739cd9ef77ff"),
                (x"ffff9ce733b5ad6b4d294a508421084a53ab5b5a4cf2e77bff"),
                (x"ffff9ce739b5ad6b5b494a108421084a53ab5a73d4f2c633ff"),
                (x"fffffcb18ccdad6b4f494a5294210842533b5a73b659ffffff"),

                -- 7_explosion_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fff39ce73967fffce739ce739ce739cb19ffffffffffffffff"),
                (x"ce739ce739cb199ce739ce739ce739ce739fffffffffffffff"),
                (x"63339cce79ce7399ce76b4f369cf39b5ad9ce58cffffffffff"),
                (x"63339cce79ce7399ce76b4f369cf39b5ad9ce58cffffffffff"),
                (x"63333b5ad39e7339e35ad4ed6b5a739ce73ce673cfffffffff"),
                (x"ce6d6b5ad6b4e769e3539ead69ced3ce7339dad6cf7fffffff"),
                (x"b5ad6b5ad6b5ad39ce76b6ad39ce73cce76b4f396319ef7fff"),
                (x"b5ad6b5ad6b5ad39ce76b6ad39ce73cce76b4f396319ef7fff"),
                (x"b5ad6b5ad6b4e694ea76b4f58c613ab5ad6b5b39ce7def7fff"),
                (x"b5ad6b4e73b6b494a756b69294a53a9eb53b5b39ce739cffff"),
                (x"9ced3d631ad25294a716b4d294a75ad2529d4e73ce739cffff"),
                (x"d6b494a5294a5294a53ad69294a538d2529d4ed69ced39e7ff"),
                (x"4a52942529c2529c61294a5384a7094e31ac6b5a9ced39e73f"),
                (x"4a52942529c2529c61294a5384a7094e31ac6b5a9ced39e73f"),
                (x"4a509421084a1094a5294a109c6129d4e7ad6a73b4ed6b5a7f"),
                (x"4a50842108421094a138c21094a529c4e7a9dad6b5ad6b5a7f"),
                (x"4a50842108421084210842108421084eb539dad6b4ed6b4f3f"),
                (x"4210842108421084210842108421294a53a9ced69ced6b659f"),
                (x"4210842108421084210842108421294a53a9ced69ced6b659f"),
                (x"4210842108421084a508421084a7094a5294ced6b5a79ce59a"),
                (x"421084a5294a108425294a5294a538d2529d4ed6b5a79ce7da"),
                (x"421294a5294a52842718c63184a538d6b49c4ed6b5b39ce733"),
                (x"4a5294a5294e309c25294a529c613ab5ada4ced6b6739ce7fa"),
                (x"4a5294a5294e309c25294a529c613ab5ada4ced6b6739ce7fa"),
                (x"9cf5a9ce7ac63184a7539e13a9cf499ce7ac4f39ce739cfff3"),
                (x"b5ad6b5ad69ce7ad6276b6b56b5b09c631a9ce73ce72c67ff3"),
                (x"b5ad6b4e73d4e739ea739eb13b5a7ad6b53b5ad6ce58e77ff3"),
                (x"9ce7a9a53ab4e79b5adad2756b5ad6b5ad6b5ad6cb3bfffff9"),
                (x"9ce7a9a53ab4e79b5adad2756b5ad6b5ad6b5ad6cb3bfffff9"),
                (x"b5b499eb539e739b5a7ad4ed6b5ad6b5ad69dad6cfbfffffff"),
                (x"ce6739e739cb1999dad6b5ad3b5ad69ce73cce739fffffffff"),
                (x"633396319963199cce79ce7399ced6b6739ce58cffffffffff"),
                (x"ffd8ef7bccce739ce73deb339ce733b6739677ffffffffffff"),
                (x"ffd8ef7bccce739ce73deb339ce733b6739677ffffffffffff"),
                (x"ffd9eeb18ccffffcb3fffb339ce739fffecf7fffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_1_2
                (x"ffffffb199b4e76b4d28421084a5294eb53b5ad6cb199cffff"),
                (x"ffffffb199b4e76b4d28421084a5294eb53b5ad6cb199cffff"),
                (x"fffec66733d4e76b69294a108421084eb56b5ad6b6739ce7ff"),
                (x"ffffe767334eb56b69294a108421094a533b5ad6b4f39ce7ff"),
                (x"ffffdf31939ce76b4d294a508421084253ab5ad6b5b39ce7ff"),
                (x"fffecf3199d2533b4d294a508421084a5389dad6b5a79ce7ff"),
                (x"fffecf3199d2533b4d294a508421084a5389dad6b5a79ce7ff"),
                (x"fffec667399eb53b69294a508421084a53a9dad6b4f39ce7ff"),
                (x"ffff9cb1999dada9e1294a50842109c253ab5ad6b4f39cb3ff"),
                (x"fffffcb18ccce739e3094a108421084a529d4ed69e72c67fff"),
                (x"fffffcb18ccce739e3094a108421084a529d4ed69e72c67fff"),
                (x"fffffce739ce733d612842108421294a5294a673b4f39cffff"),
                (x"ffff9ce733b5ad3d27084212842129c25294a6739ce79ce7ff"),
                (x"fffeccce76b5adac25294a52842109c25294ea73c6279ce7ff"),
                (x"fffffcce769dad39e938c2508421294a538d4e73d6a79ce7ff"),
                (x"fffffee736d6b53b4d38c2508423094eb56b5ad69ead9ce7ff"),
                (x"fffffee736d6b53b4d38c2508423094eb56b5ad69ead9ce7ff"),
                (x"fffec667369a53ad6138c2508421084eb53d4f5ad4e79ce7ff"),
                (x"ffff9ce736b6b58d2538c2508421084a5294ead6b5b39ce7ff"),
                (x"ffff9ce733b5ad3b6938c250842129c25294e273b5ad9ce7ff"),
                (x"ffff9cce76b5ad6b4f094a528421384a5294e2739da79ce7ff"),
                (x"ffff9cce76b5ad6b4f094a528421384a5294e2739da79ce7ff"),
                (x"ffff9cdad6b5ad3c69294a70942129c253a4a673b4f39ce7ff"),
                (x"ffff99dad6b5ada4a758c6129421294e31ad6a739cf39ce7ff"),
                (x"fffffb5ad3b5adac4edad69294a71a4eb5a9db39cced9ce7ff"),
                (x"fffffce733b5adac4edad2529d6a73c2529d5a73cced9cb3ff"),
                (x"fffffce733b5adac4edad2529d6a73c2529d5a73cced9cb3ff"),
                (x"fffecce733b5ad3d6b494a53a9cf5ad25299dad69cf39cffff"),
                (x"ffffe667399dad69e138c69339ce7ac6b5ab5ad69e73ffffff"),
                (x"fffffee733b5ad69ce739ce73b5adad4e73b5a73b673ffffff"),
                (x"ffffffb193b5ad69e6d6b5ad6b5ad3d5ad3ce739b4d9ffffff"),
                (x"ffffffb193b5ad69e6d6b5ad6b5ad3d5ad3ce739b4d9ffffff"),
                (x"fffffffff3ce739ce6d6b5ad3b5ad69ce79ce58cce7fffffff"),
                (x"fffffffffff3199ce736b5ad39ced39ce79ce58cefffffffff"),
                (x"ffffffffffff7acce739cce76b5ad6b5ad9cf98cffffffffff"),
                (x"fffffffffffffee66739ce736b5ad69ce79cfbdeffffffffff"),
                (x"fffffffffffffee66739ce736b5ad69ce79cfbdeffffffffff"),
                (x"ffffffffffffffffff39ce7399ced6ce73ffffffffffffffff"),
                (x"fffffffffffffffffff9cf98cce673cfffffffffffffffffff"),
                (x"fffffffffffe7339cf539eb5ffffffffffffffffffffffffff"),

                -- 7_explosion_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffff33fffe739ce72cfffeccffffcb19def99f"),
                (x"ffffffffffffffd66736b4f39ce72cee739ce739cb3def399f"),
                (x"fffffffffffb199ce736b5ad3ce739cce73ce58c6658c6672c"),
                (x"fffffffffffb199ce736b5ad3ce739cce73ce58c6658c6672c"),
                (x"ffffffffff9ce73cce739dad69ced6b5ad69e58cce7339ce79"),
                (x"fffffffffecdad69dad6b5ad6b5ad3d4e76b67399cf539a756"),
                (x"ce7ffff7accdad6b5ad6b5ad6b5b49d5ad6b6673b69339ea73"),
                (x"ce7ffff7accdad6b5ad6b5ad6b5b49d5ad6b6673b69339ea73"),
                (x"9cfff73199cdad6b4f5ad6a769cf1a9ce7a9ce73d4e76b5ad6"),
                (x"9cfff66739cce739eb18c2716b5b5ab4e78d6a739dad6b5ad6"),
                (x"9cfffce739ce733c6a739a753d69389eb494e318c6a739eb53"),
                (x"d6bf9ce739b5ad34ead6b69384a5294a529c27184a5294a529"),
                (x"9cf39ce736b5ad3c275ad6129c6318c6309421294a5294a528"),
                (x"9cf39ce736b5ad3c275ad6129c6318c6309421294a5294a528"),
                (x"d6bd9cce76b5ad3d253ad61294a5294a529421084a5294a108"),
                (x"d6999cce76b5ad34a5294a70942108421094a1084210842108"),
                (x"ffd99b5ad39dad39e9294a5284210842108421084210842108"),
                (x"fff33b5ad3b5ad69cf494a1084210842108421084210842109"),
                (x"fff33b5ad3b5ad69cf494a1084210842108421084210842109"),
                (x"ffe76b5ad6b5ad69ea78c25294a508c25284a5084210842109"),
                (x"ffe76b5ad3b4e7ad6a7ad25384a5084a5294a5084a10842509"),
                (x"fff399dad39eb5ac6b094a709c61294a538c2529c252842529"),
                (x"ffff99dad39dad3d253ad61294a53ad25294a5294a5294a75a"),
                (x"ffff99dad39dad3d253ad61294a53ad25294a5294a5294a75a"),
                (x"fffffce739cce73d253ad6b494a533b63094a529d6b1ad4ed3"),
                (x"fffffce739ce736b4f539e9294a53ab6b494a75ab4e76b5ad6"),
                (x"ffffff7bd9ce736b5ad6b6938c6353b4e7a4a673b5ad6b5ad6"),
                (x"ffffff318c66733b5a79cce739cedab4e739ced6b5ad6b5ad6"),
                (x"ffffff318c66733b5a79cce739cedab4e739ced6b5ad6b5ad6"),
                (x"fffffffffdcdad69cf39cced3b5ada9eb589da73b5ad6b5ad9"),
                (x"ffffffffffcce79cce739ce76b5ad3d6b589cf399ced6b4f2c"),
                (x"fffffffffffb199ce6d6b6733b5b33b4e739e739ce679ce72c"),
                (x"ffffffffffffffffe739ce739ce739ce739ce58cce739ce739"),
                (x"ffffffffffffffffe739ce739ce739ce739ce58cce739ce739"),
                (x"fffffffffffffffffd99ce739ce739ce739cffff66739ce73f"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_2_0
                (x"fffffffffffffffffffffe73e6319867bdffffffffffffffff"),
                (x"fffffffffffffffffffffe73e6319867bdffffffffffffffff"),
                (x"ffffffffffffffffffec667399ced6cb18cfffffffffffffff"),
                (x"fffffffffffffff7318c667399ced69e739cfbdeffffffffff"),
                (x"ffffffffffffffe66679ce7399ced6b5ad3cb18ccfffffffff"),
                (x"ffffffffffffbdecced6b5ad6b5ad39dad3ce739cfbfffffff"),
                (x"ffffffffffffbdecced6b5ad6b5ad39dad3ce739cfbfffffff"),
                (x"ffffffffff77bd9cdad6b4e73b5ad3c4e76b6739cb19ffffff"),
                (x"fffff9e72c76739cdad6b4ed39ce78421189dad6b598c67fff"),
                (x"ffffff319966733cdadad4edac630942118b5ad6b5a6c67bff"),
                (x"ffffff319966733cdadad4edac630942118b5ad6b5a6c67bff"),
                (x"fffffff7acf31969cf494e3584a52942109d5ad6b4f3debbdf"),
                (x"ffffffe73966736b5a694a529c612942108c4ed6b4f2c633df"),
                (x"fffff667369ce76b59294a1084a52842108d4ed6b5b39cb3df"),
                (x"fffffce736b5ad6b4d084210842108421084a75ab5a79ce59f"),
                (x"fffffcce73b5ad6b4d28425084210842108c275ab5ad39cf3f"),
                (x"fffffcce73b5ad6b4d28425084210842108c275ab5ad39cf3f"),
                (x"fffffcce799ce73b4d284212842108425294a75a9cf339e73f"),
                (x"fffffce739cce739e92842509421084a5284275ad6b59ce73f"),
                (x"ffff9ce739cdad6d2718c2508422e84252842673d6a739e73f"),
                (x"ffd99ce7399ce7ac25294a108bdc374210844ed69ced9cb3df"),
                (x"ffd99ce7399ce7ac25294a108bdc374210844ed69ced9cb3df"),
                (x"fff399e7339eb494a118c2108422e1ba1094ea739ce6c63bdf"),
                (x"fff39b5ad6b6b494a1294a11bbdee1ba1084ea739ced9cbbdf"),
                (x"fffbdcce739ce73d250842101bdd1bda1094e1294ce79cb3df"),
                (x"ffffe64e694eb53d210842101bdd08425384a1084ced9cb1df"),
                (x"ffffe64e694eb53d210842101bdd08425384a1084ced9cb1df"),
                (x"fffff6673ad6b5ad250842117ded0842108421084ce79cf7df"),
                (x"fffff66736b5ad6c210842108421084210842129d4f3debbff"),
                (x"ffffe667369eb534a108421084237b421094a3184cd8e77bff"),
                (x"fffddcdad69eb494210842108dec21ba109d635ad4f39cfbdf"),
                (x"fffddcdad69eb494210842108dec21ba109d635ad4f39cfbdf"),
                (x"fffcccce76b4e784a108422fbbdc210a109c275ad4ed9cfbdf"),
                (x"fffde66736b4e694a50842377086f70dee89ce734ced39e7df"),
                (x"fff39cdad6b4e694a508422f7bdd170ef68c6a739db39ce59f"),
                (x"ffff9ce733d4e7a4a5084237708421ba109c2718b5a79ce73f"),
                (x"ffff9ce733d4e7a4a5084237708421ba109c2718b5a79ce73f"),
                (x"ffffd67bd99dada4e10842377bdef70dee89ce73b5a79ce73f"),
                (x"ffddece733d4e7a4a7094a2f708421bef684eb5ab5a79ce59f"),
                (x"ffd9967bd99dada4e3094a37bbdc37da10842673b5a79ce5df"),

                -- 7_explosion_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"631dffe73ef7bdfffffdee72cfffffffffffffffffffffffff"),
                (x"ce7ddce73e677befffddee739ce7ffffffffffffffffffffff"),
                (x"6332cce72cce72c63199cda79ce739ce72cfffde9fffffffff"),
                (x"f7b3ecdad99dad9ce6739db39ce7339e739cf58ccfffffffff"),
                (x"f7b3ecdad99dad9ce6739db39ce7339e739cf58ccfffffffff"),
                (x"ce6799dad6b5ad6b69339da79ce7399dad6cb33967ffffffff"),
                (x"9cf53d5ad6b4e73b69339da73ce733b5ad36798c73bfffffff"),
                (x"b5a769ce739eb5ab6b539eb53b5a73b5ad3cb339cfbdffffff"),
                (x"b5a769ce739eb5ab6b539eb53b5a73b5ad3cb339cfbdffffff"),
                (x"d6b5ad2529c2533b6a739a53ab5a73b5ad6b5a73ce7def7fff"),
                (x"4a5294a5294a109c6b5ad2538d6a76b5ad6b4f39ce72c63bff"),
                (x"c61384a52942108425094a1094a7539ce76b4ed6b5a79cb3ff"),
                (x"c630842108421084210842509c61294a1099ead6b5ad39b3ff"),
                (x"4a52842108421084210842709c6108421094a75ab5ad9cb19f"),
                (x"4a52842108421084210842709c6108421094a75ab5ad9cb19f"),
                (x"42108421084210842108421084a5284a1084e2739ced9ce739"),
                (x"deefbddefbba108421084210842109421084ead6b4ed9ce739"),
                (x"deef7bdef7da10845c210ed0842128421084e35a9ced9ce73e"),
                (x"bdc370dee1bef6846ef7bdd174210842109c27189dad39ce6c"),
                (x"bdc370dee1bef6846ef7bdd174210842109c27189dad39ce6c"),
                (x"084370a1170843b4210845ee1bdd08421094a7189dad6b5acc"),
                (x"bdc370def70843b4211bd843742108421084a529c4e76b5ad8"),
                (x"deee1b84210dee84211bddee842128421084210846276b4f2c"),
                (x"4237746f774210842128421084a529421084210844ed6b659e"),
                (x"4237746f774210842128421084a529421084210844ed6b659e"),
                (x"421084a1084a529423094a128421094210842718c5a739e59f"),
                (x"42133c6313c6b49421294a52842109c253ac6ad69db39ce7ff"),
                (x"4a7534eb534e30842118c6b534a5294a5339dad6b672c67bff"),
                (x"9cf53c4e73d6b584a1094ce769cf5ad6b56b5ad6b672c67bff"),
                (x"9cf53c4e73d6b584a1094ce769cf5ad6b56b5ad6b672c67bff"),
                (x"b5ad6b4e69d6b49d25294ce73d6b53b5ad6b5ad6b6739cffff"),
                (x"b5ad6b5ad39ce739ce739ce73d6b53b5ad69ced6b33dffffff"),
                (x"9ce739e736b672ccced39da769cf59b4e79ce673633fffffff"),
                (x"ce739ce733ce72eee739ce5999cf339e7396758c67ffffffff"),
                (x"ce739ce733ce72eee739ce5999cf339e7396758c67ffffffff"),
                (x"ce739ce739f7bde7758c639ccce7399e72c63bdeffffffffff"),
                (x"73999cb19ef7bdfff9def7bdece739cb19ef7bffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_2_2
                (x"ffdd9cce76b4e694211bddc37def684e3184ead69e7cc6659f"),
                (x"ffdd9cce76b4e694211bddc37def684e3184ead69e7cc6659f"),
                (x"ffd99cce76b6b5a4a377b8421bdee84e3094ea73d4f39cf9df"),
                (x"fff39cce76b4e739a2e10def7bdf68421184ead69e7cc677ff"),
                (x"fff39cce76b6309c2517b8421bdf68421094ea73d4f39ce7ff"),
                (x"ffd99ce7369ce7ac23610dd17bdee8421094a673b5ad9ce73f"),
                (x"ffd99ce7369ce7ac23610dd17bdee8421094a673b5ad9ce73f"),
                (x"fffd99dad34ce739a2e10dee1bdf68421094a673b5b2c67bdf"),
                (x"fffdecdad3d6b49c250108437deee8421084e273b5a79cb3df"),
                (x"fffdece733d6b58d2517b843b42108421084275a9dad9cf7df"),
                (x"fffdece733d6b58d2517b843b42108421084275a9dad9cf7df"),
                (x"ffffe731934e3084a50846f6842108421084cf5a9db2c67bff"),
                (x"fffeeee733d252842108421084210842108c5ad6b5b2c67fff"),
                (x"fffddcce734a108421084211bbdd0842109d6b5ad6b2c67fff"),
                (x"ffdcccdad34a1084e128421170850842108d4f5a4a66c67bff"),
                (x"fffcccce734a5384a51bded170850842109d4e739ce79cf7bf"),
                (x"fffcccce734a5384a51bded170850842109d4e739ce79cf7bf"),
                (x"fffcecdad39ce7a4a117b86f7ded084a5284a75ab5ad6b673f"),
                (x"fffce64e739ce7a4a517b86e842108c21084a75a9cf339e73f"),
                (x"fffcccdad39dad34210845c37421084a529c6a739e739ce59f"),
                (x"fff399ce7ad4e6942128422e842109c6309d5ad6ce739ce7ff"),
                (x"fff399ce7ad4e6942128422e842109c6309d5ad6ce739ce7ff"),
                (x"fff39ceb5ad6b49421294a1084a5094253a9ce73ce739cffff"),
                (x"fff399e7339eb494a528421084212842533b4e739e679cffff"),
                (x"fff339dad6b6b49c2108421084210942533b5ad6b4e79cffff"),
                (x"ffd99cce76b6b494a108421084210842113b5ad6b5b39cffff"),
                (x"ffd99cce76b6b494a108421084210842113b5ad6b5b39cffff"),
                (x"fffccce736b5ad3d210842129421084a536b5a739db2c67fff"),
                (x"fffcc66733b5ad3c2108425384a5294ce76b5b396673ffffff"),
                (x"fffceee733b5ad6d250842529c63584eb539d98cf33bffffff"),
                (x"ffffe64e76b5ad6b610842718d6ad3d5ad6ccf396659ef7fff"),
                (x"ffffe64e76b5ad6b610842718d6ad3d5ad6ccf396659ef7fff"),
                (x"fffff63196b5ad69e108462739ced3b5ad6ce739733339ffff"),
                (x"ffffffb18cce739b5a78c4ed69ce73b5ad6ce7de77ffffffff"),
                (x"fffffffffece739cced39ced6b5ad6b5ad3cfbdeffffffffff"),
                (x"ffffffffffcb18ccced6b5ad3ce739cce7967bffffffffffff"),
                (x"ffffffffffcb18ccced6b5ad3ce739cce7967bffffffffffff"),
                (x"ffffffffffffbdece7339dad3ce7396318c77fffffffffffff"),
                (x"ffffffffffffffffb199cdad3ce73967ffffffffffffffffff"),
                (x"ffffffffffffffffffcc6618cf7b39ffffffffffffffffffff"),

                -- 7_explosion_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffef7999ce739f7bdef39defffdef7999ce58e"),
                (x"ffffffffffffbce633339e739631ce6319d77bdef6739ce739"),
                (x"ffffffffff6319d667339cf33ce599ce739ebb39ccf39ce739"),
                (x"ffffffffec64e79ce676b6753b5a769dad3cb339b5b339ce73"),
                (x"ffffffffec64e79ce676b6753b5a769dad3cb339b5b339ce73"),
                (x"fffffffbccb5ad39dad6b4f5a9ce739ce739ce739ced6b5ad6"),
                (x"fffffce739b5ad6b5ad6b4f5a9ce734a529d275ad2676b5ad6"),
                (x"ffffe66739b5ad6b5b5ad6b53b5a734a1084e35ad4e78c4f53"),
                (x"ffffe66739b5ad6b5b5ad6b53b5a734a1084e35ad4e78c4f53"),
                (x"ffffe66739b5ad69cd294a5299cf5ac2108423184cf494cf49"),
                (x"ffff9ce7369dadac6938c2508421294a5284275ac4f18c4d28"),
                (x"ffd999ce76c63094210842508421284e308425294a1094a108"),
                (x"f7999b5ad342108421084252942108425284210845f6845f68"),
                (x"63333b4e78421084210842128422f7da108422f708437b86fb"),
                (x"63333b4e78421084210842128422f7da108422f708437b86fb"),
                (x"c62d6b4e73c25294a10842108bdc21da10846c210dee10dc37"),
                (x"632d6b5ad69e3094a50842117086f74210846c210dd010dc21"),
                (x"632739dad69e309c250842108bdd17bdefb4237bb86e10dc37"),
                (x"f7b39cdad39eb584a108421284211b0843742108ddef7bdefb"),
                (x"f7b39cdad39eb584a108421284211b0843742108ddef7bdefb"),
                (x"ce739cdad3b5ada4a10842508421084210842108beefbdeefb"),
                (x"ce739cdad39ce784a1094a1294210842108421084210842108"),
                (x"ffd8ccdad6b6b494a508421184a70942108421084210842129"),
                (x"fffec9dad6b5ada9a5094a5384a50942108421084210842318"),
                (x"fffec9dad6b5ada9a5094a5384a50942108421084210842318"),
                (x"fffeccce76b5ad3b5a739cf494a5084a10942108425294e138"),
                (x"fffee66739ce733b5ad6b5a7ac6129d6b5ac25084a5294a529"),
                (x"ffffff7bd9cce76b5ad6b4e76d69299ce7ab4d29c253ad6b5a"),
                (x"fffffffbdece72ccced6b4e769cf5a9eb5ab6b5a9ce739da76"),
                (x"fffffffbdece72ccced6b4e769cf5a9eb5ab6b5a9ce739da76"),
                (x"ffffffffee7319e64ed6b4f399ce769a53ab4e73b5adad4f53"),
                (x"ffffffffff6672ccdad39e739ce6769a53ab5ad6b5ad39e679"),
                (x"ffffffffffcb19dce7339cf39ce7369ce79ce6d69e6d9cfb3e"),
                (x"ffffffffff9fbdffb339ce739ce676cb18c63339cb339cb32c"),
                (x"ffffffffff9fbdffb339ce739ce676cb18c63339cb339cb32c"),
                (x"ffffffffffffffffffffffff9ce739efbdfffbbd67b39cf7d9"),
                (x"fffffffffffffffffffffffff63339efffffffdef7b3fffdcc"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_3_0
                (x"ce7ffffffffffffee739ce6739cf334a529d7fffffffffffff"),
                (x"ce7ffffffffffffee739ce6739cf334a529d7fffffffffffff"),
                (x"fffffffffffffffce6739ced6b5b339ce7a67fffffffffffff"),
                (x"ffffffffffb5ad9cdad6b5ad6b5ad3ce739633ffffffffffff"),
                (x"fffffffff6b5ad69ced6b5ad6b5ad39ce769ce73ffffffffff"),
                (x"ffffffdad6b4e7a4ead6b4e769ced69dadad598cf7ffffffff"),
                (x"ffffffdad6b4e7a4ead6b4e769ced69dadad598cf7ffffffff"),
                (x"ffffffce7a9ce694ea76b4e76d6b5a9dad3c4ed6633fffffff"),
                (x"ffffffeb49d6b49c27094ced3c6138b5ada4ead6ce5dffffff"),
                (x"fffffb6b49c2108421294e2784a5299dada4e2739b3d6b7fff"),
                (x"fffffb6b49c2108421294e2784a5299dada4e2739b3d6b7fff"),
                (x"ffff9b6b49c2528421094e3494a508425294e129d66d6b33ff"),
                (x"ffff39e3094a5284a5084252942108421084a5299dad6b67ff"),
                (x"fffecceb494a1084a5284210942108421094a273b4f2c633ff"),
                (x"ffffecce7a4a528425284210842108421084275ab5b39cb3ff"),
                (x"ffffdcdada4a1084a508421084211b421084275ab5ad6b67ff"),
                (x"ffffdcdada4a1084a508421084211b421084275ab5ad6b67ff"),
                (x"fffde9dada4a52842108421084237b421084235ab5ad6b67bf"),
                (x"f799db5ad3c252942117bdf68422fb4210842108c6b539cd8c"),
                (x"f7b3965ad6b6b494a117b86e1086f742108421084253ad6b39"),
                (x"ce7399ce76b6b4842117b86f7bdc3742108421084253ad4f39"),
                (x"ce7399ce76b6b4842117b86f7bdc3742108421084253ad4f39"),
                (x"ce59ef6739b6b48423610dc37def61da10842108427139cf39"),
                (x"ffd8ef3199b4e6846c210def708517ba1084a1084ea6c6333f"),
                (x"ffffef31934a52846ef7ba11708421da1094a5294cedef3bff"),
                (x"ffffe6672942109c236846ef708421da108421084cecc67bff"),
                (x"ffffe6672942109c236846ef708421da108421084cecc67bff"),
                (x"fffeeece78421094a117bdee1086e1da10842108462739fbdf"),
                (x"fffeccce684210846f77b8421bdee10dee84210842756b658c"),
                (x"ffff6b4e69421084236108437def6845ef7da10842356b4f39"),
                (x"ffff6b5ada4210842117bdef7086e8b84210ed0842356b4f39"),
                (x"ffff6b5ada4210842117bdef7086e8b84210ed0842356b4f39"),
                (x"739969ce7a4a1084251bddee108437b843b42108422739b3de"),
                (x"633d3d63094252942517b8421086fbba10842108426d9cfbdf"),
                (x"ce5999a5384252946137bdc2108437da1084210842279cfbff"),
                (x"ce7399eb534a109c251bda2e1084210ef68421294a66c63bff"),
                (x"ce7399eb534a109c251bda2e1084210ef68421294a66c63bff"),
                (x"ce7339dad34a1084a108422e108421ba10842108d4e6c67bff"),
                (x"fff33b4e784a1084210842377084210dee842108d5acc63bff"),
                (x"ffffa9eb49d21084210842117bdc21ba108421089dacc63bff"),

                -- 7_explosion_3_1
                (x"ffff9ce72c77fffffffffff39f7bdffffffffffffffffffff9"),
                (x"ffff9ce72c77fffffffffff39f7bdffffffffffffffffffff9"),
                (x"fff39cb19e67fffffffffb199ce59effffffffffffffffffff"),
                (x"d6a73ce733b5ad663bdef3bd9ce7beefbcc9e7ffffffffffff"),
                (x"9ced39ce7a9dad6cf59ef7bd3632d3ce7399dad6ffffffffff"),
                (x"d6a76d25389dad39cf2c63333b5ad6b4e7ac6b5ad4edffffff"),
                (x"d6a76d25389dad39cf2c63333b5ad6b4e7ac6b5ad4edffffff"),
                (x"4a7139e309d6b49461339e736b5a7ad6b494a5294ead6b7fff"),
                (x"d69294a1084a108421094dad6b5b094a5294e318d4ed6b5bff"),
                (x"421084252942108421094cf5ad6929425284a508d4e76b5bff"),
                (x"421084252942108421094cf5ad6929425284a508d4e76b5bff"),
                (x"421084a5294210842528421084a52842108421084a756b67ff"),
                (x"42109c21084210842708421084a5084a1094a108c25339e73d"),
                (x"421084e3094a108da11bded08421084a5294a1084eb539db39"),
                (x"42108425284211bda377b8768421084252942129c4ed6b5a79"),
                (x"42108ddef7ddee1bdd17b8437bdee842108425294dad6b5a79"),
                (x"42108ddef7ddee1bdd17b8437bdee842108425294dad6b5a79"),
                (x"4210845ee1bdee10df6845ee1086e8421084e3189ce76b5a79"),
                (x"42377b8421bdee10dee845c37bdf68421084ea73b4e76b5ad3"),
                (x"bdee1084210def7086f7bdef708508421094a7189dad6b5ad3"),
                (x"bdc21084210843bb842108777085084210842529c6a76b5ad3"),
                (x"bdc21084210843bb842108777085084210842529c6a76b5ad3"),
                (x"08421084370defbbdc210a361bdefb42108421294ead6b5b39"),
                (x"084210defbba108084210dc37bdf7bda10842129c6ad39ce73"),
                (x"bdc370ef77bdee80ef7bddf68421084210842273b4e739e669"),
                (x"422e8da10808437ba108421084210842108426d6b5ad39e669"),
                (x"422e8da10808437ba108421084210842108426d6b5ad39e669"),
                (x"4210842108d8437421094a10842108421094275ad4f56b6749"),
                (x"42108421084043b421094a50842108421094a5294e3539b19a"),
                (x"421084210846f68421094a108421084a5284e318d4ed39b3ff"),
                (x"421084a10842108421094a1084211ad6b534a673b59939ffff"),
                (x"421084a10842108421094a1084211ad6b534a673b59939ffff"),
                (x"9cf5a4a10842108421294a50842316b5ad69ea73cb3dffffff"),
                (x"b5ad34a109421084e2739e9294a756b5ad3b658ccb3fffffff"),
                (x"b5ad39ce769eb5ad4ed6b4f094a756b6739b5bde77ffffffff"),
                (x"6318c667399dad6b4d9ef327ad6a76b672cb5ad6ffffffffff"),
                (x"6318c667399dad6b4d9ef327ad6a76b672cb5ad6ffffffffff"),
                (x"739de77bde64e73cfbce73273d6a79cb18ccb3ffffffffffff"),
                (x"fffffffffef673967bfffe739ce59dffffffffffffffffffff"),
                (x"fffffffffff673967ffffff39ce59fffffffffffffffffffff"),

                -- 7_explosion_3_2
                (x"fffee65ad69a10842117b8437bdd084210842108d27539ebff"),
                (x"fffee65ad69a10842117b8437bdd084210842108d27539ebff"),
                (x"fffee65ad6d2108422e108421bdf6842108421084e276b4f3f"),
                (x"ffffe64e73d210842117b8421086e8421084a1084ced39cf39"),
                (x"fffee64e694a5284236108421086e8da109c25084cf539e739"),
                (x"ffffecce68421084211bddc2108437ba53842529461339e599"),
                (x"ffffecce68421084211bddc2108437ba53842529461339e599"),
                (x"fffdecdac94210842117beee108421ba109425294271ad4fcc"),
                (x"f7bcc9ce684210846c37bdc21086f7da109421084ea739d98e"),
                (x"ce733b6b484211b08437ba2e1bdef7ba1084210846ad6b5bff"),
                (x"ce733b6b484211b08437ba2e1bdef7ba1084210846ad6b5bff"),
                (x"ce733b6b4842108ddee84237bbdc210ef684210842676b5bff"),
                (x"63199b6b4942108422e1086f708421bef7b4210842279cb3ff"),
                (x"fffde9ce78421084211bd86e1086f7ba1084a5084627debbff"),
                (x"ffffe65ad34a1084211bd8421bdefb46f68c25084272c67bff"),
                (x"fffeef5ad34a5294a51bd8421bdd08bdefb421294cd9ef7bff"),
                (x"fffeef5ad34a5294a51bd8421bdd08bdefb421294cd9ef7bff"),
                (x"fff2c64e7a4a1084a117bdd01bdef70843b42273b659ef399f"),
                (x"ce7339e309421084211bd877bbdc370ef684235ab673ef7999"),
                (x"ce733d2529421084210845c37bdee1ba1084235ab5a739e739"),
                (x"ce73ad2529421084210845ee1086e1ba1084a75ab5acc6673e"),
                (x"ce73ad2529421084210845ee1086e1ba1084a75ab5acc6673e"),
                (x"631939eb5ac21084210846ee842377ba10842529c4ed6b759e"),
                (x"fffb9b5ad6b6b484210846f684210842108421294ead39fbdf"),
                (x"ffff9b5ad6b6b494210846d0842108421094a1084ead9cf7ff"),
                (x"fffecce736b6b4942108421084210842529421294ea79cfbff"),
                (x"fffecce736b6b4942108421084210842529421294ea79cfbff"),
                (x"fffec66733b4e684a508421084a508425294a1084a759cb3ff"),
                (x"ffff9b5ad69a5294a108421084a529421094a1294a7139cfff"),
                (x"fffecb5ad9d25384a528421094a7584a10842129c2756b67ff"),
                (x"fffffb7bcc9ce784ead39a529c62784a52842108c2756b7fff"),
                (x"fffffb7bcc9ce784ead39a529c62784a52842108c2756b7fff"),
                (x"ffffffb9d9cdada4ead6b61389ced34e309c275ad275ffffff"),
                (x"ffffffffec65ad3c4ed39eb5ab5a73b4e7a4a6739ea7ffffff"),
                (x"fffffffffff3196d6ad39dad3b5a73b5ada4ea73b5adffffff"),
                (x"fffffffffffce739da739ced6b5ad6b5ad39dad6b5bfffffff"),
                (x"fffffffffffce739da739ced6b5ad6b5ad39dad6b5bfffffff"),
                (x"fffffffffffffec66739cced6b5ad6b5ad6ce6d6b7ffffffff"),
                (x"fffffffffffffff66a739cf36b5ad39ce79cffffffffffffff"),
                (x"fffffffffffffffd25294cf339ce79ce739efffffffffffff9"),

                -- 7_explosion_3_3
                (x"ffffffffffffffffffffffd99ce73ffffff66739f7ffffffff"),
                (x"ffffffffffffffffffffffd99ce73ffffff66739f7ffffffff"),
                (x"ffffffffffffffffffffff599ce739ffffe66739f7bfffffff"),
                (x"fffffffffffffeccb199ce67a9ce6c77bdecce7367bce779ce"),
                (x"fffffffffffdad6b3336b5a7ad6a6cf3193b5ad69e72c6318c"),
                (x"ffffffffff77bd6b6736b5b494a713b5ad3d6b5a9da739ced6"),
                (x"ffffffffff77bd6b6736b5b494a713b5ad3d6b5a9da739ced6"),
                (x"ffffffffeccb199b4ed6b5b494a53a9ce784a108425094ced6"),
                (x"fffffffbcccce7a9dad6b5b08421094a52842108421094eb53"),
                (x"fffff9b196b4e694cf5ad6908421084a10842108421094a108"),
                (x"fffff9b196b4e694cf5ad6908421084a10842108421094a108"),
                (x"fffec9dad3d63184a1294a108421084a1084237b4210842108"),
                (x"d698c9eb584a5294a50842108421094a10846c214210842108"),
                (x"4a759b6b53d6b494250842108421084a10845c21da10842108"),
                (x"4a6799dad6b5ac942108421084210842108bdc210a11bda2e8"),
                (x"4a6799ce73b4e68421084210842377def7b0a2f7bdf610dc37"),
                (x"4a6799ce73b4e68421084210842377def7b0a2f7bdf610dc37"),
                (x"9ce739dadac25284211bdef77bdc37084210a108beee108421"),
                (x"ce736b5ada4a5284210846ef70876808437beef70dc2108421"),
                (x"9ced6b4e7ac25294210842101bdf6108421bec210842108437"),
                (x"9ced6b5ad69e3094a50842101bdef7bdee10def708421086f7"),
                (x"9ced6b5ad69e3094a50842101bdef7bdee10def708421086f7"),
                (x"9ced6b4e73b4e7a4a10842377bdc3745ef7086f7b8437bdf68"),
                (x"ce676b4e739e3184a108422e1086f746f77086f7b86e842108"),
                (x"ce676b5ad64a52942108422f7bdc21ba117b86f7ddefbda108"),
                (x"ce676b5ad3c2528425284210842361bef68ded084212842108"),
                (x"ce676b5ad3c2528425284210842361bef68ded084212842108"),
                (x"ce7369eb5a4a1084a5294a1084211bda108da1084a7094a108"),
                (x"ef7399a529c21084a5094a10942108463094210842118c2508"),
                (x"ffff9b6b494a1084210842129421084252942108425294a108"),
                (x"ffff6b4e73d21094a1284253ad6b534a108421084252842108"),
                (x"ffff6b4e73d21094a1284253ad6b534a108421084252842108"),
                (x"ffff6b5ad3d63184a5294a716b5ad64a108421084a1094a53a"),
                (x"fffffb5ada4a5294a75ad6a76b5b399a5384275ad27139cf09"),
                (x"ffffffdad3d6b5ac6a76b5ad69cf2c667339ced69e13ad5a7a"),
                (x"fffffffffffdad69e739ccecc9cfdef319dcdad69ea739ced3"),
                (x"fffffffffffdad69e739ccecc9cfdef319dcdad69ea739ced3"),
                (x"ffffffffffffff99b3ddefbb9ce7cef7bce65ad6b4f39cce7a"),
                (x"ffffffffffffffffffffff999ce58cffffffffff67999ce73f"),
                (x"ce7ffffffffffffffffffffdece73fffffffffff73339ce7ff"),

                -- 8_bonus-life
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6f39ce739ce71ad6b5bce739ce739c6b5ad9cca5"),
                (x"294b39b5ad6f39ce739ce71ad6b5bce739ce739c6b5ad9cca5"),
                (x"294b39b5b4a4e73c63189ce94a52939a53ad4e73a51ad9cca5"),
                (x"294b39b5b4a4e73c63189ce94a52939a53ad4e73a51ad9cca5"),
                (x"294b39b5b4a4e73c63189ce94a52939a53ad4e73a51ad9cca5"),
                (x"294b9cd2939a529421084a6739ce694a11ef6b5a9ce94ce4a5"),
                (x"294b9cd2939a529421084a6739ce694a11ef6b5a9ce94ce4a5"),
                (x"294b9cd28948421085084235ac6308439cb5fbded6a94ce4a5"),
                (x"294b9cd28948421085084235ac6308439cb5fbded6a94ce4a5"),
                (x"294b9cd2894842108508a53bda529de908e721084a694ce4a5"),
                (x"294b9cd2894842108508a53bda529de908e721084a694ce4a5"),
                (x"294b9cd2894a10842294a508484200077a8421084a694ce4a5"),
                (x"294b9cd2894a10842294a508484200077a8421084a694ce4a5"),
                (x"294b9cd2939a108bde9439ca57bdfded288421089ce94ce4a5"),
                (x"294b9cd2939a108bde9439ca57bdfded288421089ce94ce4a5"),
                (x"294b9cd2939a108bde9439ca57bdfded288421089ce94ce4a5"),
                (x"294b39b5b4a25294239c319ef739ddef38842529a51ad9cca5"),
                (x"294b39b5b4a25294239c319ef739ddef38842529a51ad9cca5"),
                (x"294b39b5bce4e73c6294003bdef7bce5298c4e73e71ad9cca5"),
                (x"294b39b5bce4e73c6294003bdef7bce5298c4e73e71ad9cca5"),
                (x"294b39b5ad6d2949cf5aa539ce7394a6b539d2946b5ad9cca5"),
                (x"294b39b5ad6d2949cf5aa539ce7394a6b539d2946b5ad9cca5"),
                (x"294b39b5ad6b5ada5294d69084211ad5294a35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ada5294d69084211ad5294a35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ada5294d69084211ad5294a35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b5adef5294a53deb5ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b5adef5294a53deb5ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b5ad6b694a528d6b5ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b5ad6b694a528d6b5ad6b5ad6b5ad9cca5"),
                (x"294b39ce739ce739ce739cf39ce7339ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739cf39ce7339ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 9_bonus-godmod
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce739ce739ce739cfbdef7b39ce79cce739ce739cca5"),
                (x"294b39ce739ce739ce739cfbdef7b39ce79cce739ce739cca5"),
                (x"294b39b5ad6b5adef694a516b21094a529deb5ad6b5ad9cca5"),
                (x"294b39b5ad6b5adef694a516b21094a529deb5ad6b5ad9cca5"),
                (x"294b39b5ad6f39c5ac841094a5ad6212d64277bd6b5ad9cca5"),
                (x"294b39b5ad6f39c5ac841094a5ad6212d64277bd6b5ad9cca5"),
                (x"294b39b5ad6d2945296ba50c65ad663294b5d2946b5ad9cca5"),
                (x"294b39b5ad6d2945296ba50c65ad663294b5d2946b5ad9cca5"),
                (x"294b39b5ad6d2945296ba50c65ad663294b5d2946b5ad9cca5"),
                (x"294b39b5ad6f39c39d4a3194a5ad74a1ceb588426b5ad9cca5"),
                (x"294b39b5ad6f39c39d4a3194a5ad74a1ceb588426b5ad9cca5"),
                (x"294b39b5ad6d2945294aa514a52954a462b5f7bd6b5ad9cca5"),
                (x"294b39b5ad6d2945294aa514a52954a462b5f7bd6b5ad9cca5"),
                (x"294b39b5bded294a539c10842318d4a5294a77bd6b5ad9cca5"),
                (x"294b39b5bded294a539c10842318d4a5294a77bd6b5ad9cca5"),
                (x"294b39d28b58421ef79c5294a8c6273c634a77bd6b5ad9cca5"),
                (x"294b39d28b58421ef79c5294a8c6273c634a77bd6b5ad9cca5"),
                (x"294b39d28a52d6b5afbd39d4a39ceb5ad6a5739c6b5ad9cca5"),
                (x"294b39d28a52d6b5afbd39d4a39ceb5ad6a5739c6b5ad9cca5"),
                (x"294b39d28a52d6b5afbd39d4a39ceb5ad6a5739c6b5ad9cca5"),
                (x"294b39d29ce294a7bd6b5adcea528a52d6b5f39c6b5ad9cca5"),
                (x"294b39d29ce294a7bd6b5adcea528a52d6b5f39c6b5ad9cca5"),
                (x"294b39b5bce18c652a520856ba528a52d718d2946b5ad9cca5"),
                (x"294b39b5bce18c652a520856ba528a52d718d2946b5ad9cca5"),
                (x"294b39b5ad6f39c3194a5ad6b1084a529463739c6b5ad9cca5"),
                (x"294b39b5ad6f39c3194a5ad6b1084a529463739c6b5ad9cca5"),
                (x"294b39b5ad6b5ade70c65296ba528a5295ce35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ade70c65296ba528a5295ce35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ade70c65296ba528a5295ce35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b69439d4a318def18cd6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b69439d4a318def18cd6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ade73bd5294a5ad6b5c63ce35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ade73bd5294a5ad6b5c63ce35ad6b5ad9cca5"),
                (x"294b39ce739ce73a539c3184210846318d4a4e739ce739cca5"),
                (x"294b39ce739ce73a539c3184210846318d4a4e739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 10_bonus-wallhack
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39e739cce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39e739cce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294a10842422d6b5af9ce73bde739ce739ce77bde739c9cca5"),
                (x"294a10842422d6b5af9ce73bde739ce739ce77bde739c9cca5"),
                (x"294b39b5ad6fbde1098c18ef718c74a31831def718e94ce4a5"),
                (x"294b39b5ad6fbde1098c18ef718c74a31831def718e94ce4a5"),
                (x"294b39b5ad6fbde1098c18ef718c74a31831def718e94ce4a5"),
                (x"294b9cb5a422d6b8416b5ac6318c74a318318c6318e94ce4a5"),
                (x"294b9cb5a422d6b8416b5ac6318c74a318318c6318e94ce4a5"),
                (x"294b39b5ad6fbde3198c6318c63194a318c6318c632949cca5"),
                (x"294b39b5ad6fbde3198c6318c63194a318c6318c632949cca5"),
                (x"294b399084214a52961000000a5294a5294a5294a52949cca5"),
                (x"294b399084214a52961000000a5294a5294a5294a52949cca5"),
                (x"294b39b5ad6fbde318c61098c18c77b8c74a0c6329694ce4a5"),
                (x"294b39b5ad6fbde318c61098c18c77b8c74a0c6329694ce4a5"),
                (x"294a109084214a55ad6b5ad6b18c6318c74a0c6318e94ce4a5"),
                (x"294a109084214a55ad6b5ad6b18c6318c74a0c6318e94ce4a5"),
                (x"294a109084214a55ad6b5ad6b18c6318c74a0c6318e94ce4a5"),
                (x"294b39b5ad6fbde6318c1098c6318c63194a318c632949cca5"),
                (x"294b39b5ad6fbde6318c1098c6318c63194a318c632949cca5"),
                (x"294b3990842421000000a5294a5294a5294a5294a52949cca5"),
                (x"294b3990842421000000a5294a5294a5294a5294a52949cca5"),
                (x"294b39b5ad6fbde6306318ef718c74a31831def718e949cca5"),
                (x"294b39b5ad6fbde6306318ef718c74a31831def718e949cca5"),
                (x"294a10908422d6b5ad6b18c6318c74a318318c6318e94ce4a5"),
                (x"294a10908422d6b5ad6b18c6318c74a318318c6318e94ce4a5"),
                (x"294a10908422d6b5ad6b18c6318c74a318318c6318e94ce4a5"),
                (x"294b39b5ad6ffff318c6e739ce739ce739ce739ce739c9cca5"),
                (x"294b39b5ad6ffff318c6e739ce739ce739ce739ce739c9cca5"),
                (x"294b9cb5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294b9cb5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 11_bonus-speed
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39b5ad6b5ad6b5ada518c6318c6318c6318ce71ad9cca5"),
                (x"294b39b5ad6b5ad6b5ada518c6318c6318c6318ce71ad9cca5"),
                (x"294b39b5ad6b5ad6b5ade70630842b5c20a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b5ade70630842b5c20a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b7bd421084a53ad420a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b7bd421084a53ad420a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b7bd421084a53ad420a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b5adef6318c6318c20a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b5adef6318c6318c20a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b79c4a508c63139c20a518c6e71ad9cca5"),
                (x"294b39b5ad6b5ad6b79c4a508c63139c20a518c6e71ad9cca5"),
                (x"294b39b5ad6f39ca5294ef6318c6318c20a577bde71ad9cca5"),
                (x"294b39b5ad6f39ca5294ef6318c6318c20a577bde71ad9cca5"),
                (x"294b39b5bce77bd5ac212116b5ad6b5c20a518c6e71ad9cca5"),
                (x"294b39b5bce77bd5ac212116b5ad6b5c20a518c6e71ad9cca5"),
                (x"294b39d28632d6b0856b5ad6b5ad708294a5294affe949cca5"),
                (x"294b39d28632d6b0856b5ad6b5ad708294a5294affe949cca5"),
                (x"294b39d28632d6b0856b5ad6b5ad708294a5294affe949cca5"),
                (x"294b39d28a52d6bef694842105294a577b4a18c6ffe949cca5"),
                (x"294b39d28a52d6bef694842105294a577b4a18c6ffe949cca5"),
                (x"294b39d286377bd42108e73bd318ddea1084739ce72949cca5"),
                (x"294b39d286377bd42108e73bd318ddea1084739ce72949cca5"),
                (x"294b39b5bce21087bdce42294a528843dee72108a52949cca5"),
                (x"294b39b5bce21087bdce42294a528843dee72108a52949cca5"),
                (x"294b39b5bdea10873bdec6294e7388439def6318e71ad9cca5"),
                (x"294b39b5bdea10873bdec6294e7388439def6318e71ad9cca5"),
                (x"294b39b5bdea10873bdec6294e7388439def6318e71ad9cca5"),
                (x"294b39b5ad6f7bd42318e71ad6b5bdea118c739c6b5ad9cca5"),
                (x"294b39b5ad6f7bd42318e71ad6b5bdea118c739c6b5ad9cca5"),
                (x"294b39b5ad6b5ada52946b5ad6b5ad6d294a35ad6b5ad9cca5"),
                (x"294b39b5ad6b5ada52946b5ad6b5ad6d294a35ad6b5ad9cca5"),
                (x"294b39ce739ce73ce7399ce739ce739e739cce739ce739cca5"),
                (x"294b39ce739ce73ce7399ce739ce739e739cce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 12_bonus-addbomb
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce739ce739ce739ce739ce739ce739e739ce6739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739e739ce6739cca5"),
                (x"294b39b5ad6b5ad6b694a5294a5294a739fff7bda51ad9cca5"),
                (x"294b39b5ad6b5ad6b694a5294a5294a739fff7bda51ad9cca5"),
                (x"294b39b5ad6f39ce739cef79ce738f7f7ae710849ce94ce4a5"),
                (x"294b39b5ad6f39ce739cef79ce738f7f7ae710849ce94ce4a5"),
                (x"294b39b5bce0000ef5ef7bf9c294a4277a4214a5e71ad9cca5"),
                (x"294b39b5bce0000ef5ef7bf9c294a4277a4214a5e71ad9cca5"),
                (x"294b39b5bce0000ef5ef7bf9c294a4277a4214a5e71ad9cca5"),
                (x"294b39b5bce77bd5ac21842940842b58854a5294e71ad9cca5"),
                (x"294b39b5bce77bd5ac21842940842b58854a5294e71ad9cca5"),
                (x"294b39d29debdef08484842948421083dfce739ce72949cca5"),
                (x"294b39d29debdef08484842948421083dfce739ce72949cca5"),
                (x"294b39d28f7c2105ae107bfbda528f7b9dded294e72949cca5"),
                (x"294b39d28f7c2105ae107bfbda528f7b9dded294e72949cca5"),
                (x"294b39d28f7c210841ef7bdefef7b4a5294a5294e72949cca5"),
                (x"294b39d28f7c210841ef7bdefef7b4a5294a5294e72949cca5"),
                (x"294b39d28f7bdef7bdef7bdef7bdfdef7bded294e72949cca5"),
                (x"294b39d28f7bdef7bdef7bdef7bdfdef7bded294e72949cca5"),
                (x"294b39d28f7bdef7bdef7bdef7bdfdef7bded294e72949cca5"),
                (x"294b39d28633def7bdef7bdef739ddef7b4a5294e72949cca5"),
                (x"294b39d28633def7bdef7bdef739ddef7b4a5294e72949cca5"),
                (x"294b39d29ce77bd7bdef7bdceef7ae777b4a5294e72949cca5"),
                (x"294b39d29ce77bd7bdef7bdceef7ae777b4a5294e72949cca5"),
                (x"294b39b5bce5294ef5ce73bbdef7bded294a5294e71ad9cca5"),
                (x"294b39b5bce5294ef5ce73bbdef7bded294a5294e71ad9cca5"),
                (x"294b39b5bce0000a53bdef7bda5294a5294a5294e71ad9cca5"),
                (x"294b39b5bce0000a53bdef7bda5294a5294a5294e71ad9cca5"),
                (x"294b39b5bce0000a53bdef7bda5294a5294a5294e71ad9cca5"),
                (x"294b39b5ad6f39ce739ce739ce739ce739ce739c6b5ad9cca5"),
                (x"294b39b5ad6f39ce739ce739ce739ce739ce739c6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b694a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b694a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 13_bonus-power
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39b5ad6b5ad6b5ad6b58c6b5ad6b18d6b5ad631ad9cca5"),
                (x"294b39b5ad6b5ad6b5ad6b58c6b5ad6b18d6b5ad631ad9cca5"),
                (x"294b39b5ad6b5ad6b5ad6335a6318c6210c6318cc618c9cca5"),
                (x"294b39b5ad6b5ad6b5ad6335a6318c6210c6318cc618c9cca5"),
                (x"294b39b5ad6b5ad6318c4a508631884210c621084a7399cca5"),
                (x"294b39b5ad6b5ad6318c4a508631884210c621084a7399cca5"),
                (x"294b39b5ad6b5ad6318c4a508631884210c621084a7399cca5"),
                (x"294b39b5ad6b18cc6021085084210842108421084a58c9cca5"),
                (x"294b39b5ad6b18cc6021085084210842108421084a58c9cca5"),
                (x"294b39b5ac6631808421421080842842108421084a58c9cca5"),
                (x"294b39b5ac6631808421421080842842108421084a58c9cca5"),
                (x"294b39b5ac65ef7423bdbdd08ef7a422108421084a58c9cca5"),
                (x"294b39b5ac65ef7423bdbdd08ef7a422108421084a58c9cca5"),
                (x"294b39b1894a1084229408508a528422108421084a58c9cca5"),
                (x"294b39b1894a1084229408508a528422108421084a58c9cca5"),
                (x"294b39b18842108423de08508ef7a10a108421084a7399cca5"),
                (x"294b39b18842108423de08508ef7a10a108421084a7399cca5"),
                (x"294b39b18842108423de08508ef7a10a108421084a7399cca5"),
                (x"294b39b1884210821108421084210842108421084a58c9cca5"),
                (x"294b39b1884210821108421084210842108421084a58c9cca5"),
                (x"294b39e7294a10863294a5294a5294a210842529631ad9cca5"),
                (x"294b39e7294a10863294a5294a5294a210842529631ad9cca5"),
                (x"294b39b198c21084218cce739a5298c210846b5a631ad9cca5"),
                (x"294b39b198c21084218cce739a5298c210846b5a631ad9cca5"),
                (x"294b39b5ac66b5a421086318c4a5284211ad318c6b5ad9cca5"),
                (x"294b39b5ac66b5a421086318c4a5284211ad318c6b5ad9cca5"),
                (x"294b39b5ac66b5a421086318c4a5284211ad318c6b5ad9cca5"),
                (x"294b39b5ad6b18c6310842108421094b18c635ad6b5ad9cca5"),
                (x"294b39b5ad6b18c6310842108421094b18c635ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b58c6318c6318c635ad6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b58c6318c6318c635ad6b5ad6b5ad9cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 14_malus-inversed-commands
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739bdef7bdef7bdef7bdef9ce739ce739ce65"),
                (x"296739ce739ce739bdef7bdef7bdef7bdef9ce739ce739ce65"),
                (x"296736b5ad6bdef7ad6b5ad6b5ad6b5ad6b7bdef6b5ad6ce65"),
                (x"296736b5ad6bdef7ad6b5ad6b5ad6b5ad6b7bdef6b5ad6ce65"),
                (x"296736b5ef7ad6b5ad6b5ad6b5ad6b5ad6b5ad6b7bded6ce65"),
                (x"296736b5ef7ad6b5ad6b5ad6b5ad6b5ad6b5ad6b7bded6ce65"),
                (x"296736b5ef7ad6b5ad6b5ad6b5ad6b5ad6b5ad6b7bded6ce65"),
                (x"296737bd6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6f7ce65"),
                (x"296737bd6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6f7ce65"),
                (x"296737bd6b5bdef7ad6b5ad6b5ad6b5ad6b7bdef5ad6f7ce65"),
                (x"296737bd6b5bdef7ad6b5ad6b5ad6b5ad6b7bdef5ad6f7ce65"),
                (x"295ef5adef7bdef7bdef5ad6b5ad6b5bdef7bdef7bdeb5bde5"),
                (x"295ef5adef7bdef7bdef5ad6b5ad6b5bdef7bdef7bdeb5bde5"),
                (x"295ef5adef7bdef7bdef5ad6b5ad6b5bdef7bdef7bdeb5bde5"),
                (x"295ef5adef7ad6f7bdef7bd6b5ad6f7bdef7bd6b7bdeb5bde5"),
                (x"295ef5adef7ad6f7bdef7bd6b5ad6f7bdef7bd6b7bdeb5bde5"),
                (x"295ef5adef7bdef7d2947be94a528f7d2947bdef7bdeb5bde5"),
                (x"295ef5adef7bdef7d2947be94a528f7d2947bdef7bdeb5bde5"),
                (x"295ef5adef7bdef7d2947be94a528f7d2947bdef7bdeb5bde5"),
                (x"295ef5ad6b5bdef7d2945ae94a528b5d2947bdef5ad6b5bde5"),
                (x"295ef5ad6b5bdef7d2945ae94a528b5d2947bdef5ad6b5bde5"),
                (x"295ef5ad6b5ad6b5d294a5294a5294a52945ad6b5ad6b5bde5"),
                (x"295ef5ad6b5ad6b5d294a5294a5294a52945ad6b5ad6b5bde5"),
                (x"296737bd6b5ad6b5ad6b5ae94a528b5ad6b5ad6b5ad6f7ce65"),
                (x"296737bd6b5ad6b5ad6b5ae94a528b5ad6b5ad6b5ad6f7ce65"),
                (x"296737bd6b5ad6b5ad6b5ae94a528b5ad6b5ad6b5ad6f7ce65"),
                (x"296736b5ef7bdeb5ad6b5ae94a528b5ad6b5adef7bded6ce65"),
                (x"296736b5ef7bdeb5ad6b5ae94a528b5ad6b5adef7bded6ce65"),
                (x"296736b5ad6bdeb5d294a5294a5294a52945adef6b5ad6ce65"),
                (x"296736b5ad6bdeb5d294a5294a5294a52945adef6b5ad6ce65"),
                (x"296736b5ad6bdeb5d2945adef7bdeb5d2945adef6b5ad6ce65"),
                (x"296736b5ad6bdeb5d2945adef7bdeb5d2945adef6b5ad6ce65"),
                (x"296736b5ad6bdeb5d2945adef7bdeb5d2945adef6b5ad6ce65"),
                (x"296736b5ad6bdf4a52947bdef7bdef7d294a51ef6b5ad6ce65"),
                (x"296736b5ad6bdf4a52947bdef7bdef7d294a51ef6b5ad6ce65"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739ce65"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739ce65"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 15_malus-disable-bombs
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce79ce7399ce73ce694a5299cce739e739ce6739cca5"),
                (x"294b39ce79ce7399ce73ce694a5299cce739e739ce6739cca5"),
                (x"294b9cd294a5294ef694a510818c74a529ded294a5294ce4a5"),
                (x"294b9cd294a5294ef694a510818c74a529ded294a5294ce4a5"),
                (x"294b9cd28840c63e70e739c214211de8014a0c6342294ce4a5"),
                (x"294b9cd28840c63e70e739c214211de8014a0c6342294ce4a5"),
                (x"294b39d28319ce7843bd18c21421031d280077bd18e949cca5"),
                (x"294b39d28319ce7843bd18c21421031d280077bd18e949cca5"),
                (x"294b39d28319ce7843bd18c21421031d280077bd18e949cca5"),
                (x"294b39f39ce2d6b5ae9418d08421031d29ded294e73bd9cca5"),
                (x"294b39f39ce2d6b5ae9418d08421031d29ded294e73bd9cca5"),
                (x"294b39d29ffad6b0861018d08421031d29ded294002949cca5"),
                (x"294b39d29ffad6b0861018d08421031d29ded294002949cca5"),
                (x"294b39d29082d6b084217be94a529ef39dded294e72949cca5"),
                (x"294b39d29082d6b084217be94a529ef39dded294e72949cca5"),
                (x"294b39d29083def7bd6b5ae108420f7f7bce5294002949cca5"),
                (x"294b39d29083def7bd6b5ae108420f7f7bce5294002949cca5"),
                (x"294b39d28e70c63a51ef842107bdee75294a0c63a52949cca5"),
                (x"294b39d28e70c63a51ef842107bdee75294a0c63a52949cca5"),
                (x"294b39d28e70c63a51ef842107bdee75294a0c63a52949cca5"),
                (x"294b9cd28318421422947bdef739dce52884042118e94ce4a5"),
                (x"294b9cd28318421422947bdef739dce52884042118e94ce4a5"),
                (x"294b9cd2810842142294ef7bdef7b4a52884042108694ce4a5"),
                (x"294b9cd2810842142294ef7bdef7b4a52884042108694ce4a5"),
                (x"294b9cd28840c6318e94a5294a5294a528318c6342294ce4a5"),
                (x"294b9cd28840c6318e94a5294a5294a528318c6342294ce4a5"),
                (x"294b39b5bce0000a5294a5294a5294a5294a0000e71ad9cca5"),
                (x"294b39b5bce0000a5294a5294a5294a5294a0000e71ad9cca5"),
                (x"294b39b5bce0000a5294a5294a5294a5294a0000e71ad9cca5"),
                (x"294b39b5ad6f39ce739ce739ce739ce739ce739c6b5ad9cca5"),
                (x"294b39b5ad6f39ce739ce739ce739ce739ce739c6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b694a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"294b39b5ad6b5ad6b694a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 16_malus-remove-power
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739b5ad6b5ad6b58c6b5ad6b18c64e739ce739cca5"),
                (x"294b39ce739b5ad6b5ad6b58c6b5ad6b18c64e739ce739cca5"),
                (x"294b39ce739ce736b5ad6335a6318c663139ce739ce739cca5"),
                (x"294b39ce739ce736b5ad6335a6318c663139ce739ce739cca5"),
                (x"294b39ce739ce739cd8c4a508631894ce739ce739cf399cca5"),
                (x"294b39ce739ce739cd8c4a508631894ce739ce739cf399cca5"),
                (x"294b39ce739ce739cd8c4a508631894ce739ce739cf399cca5"),
                (x"294b39fbd39ce739ce73bdd084a5339ce739ce734a58c9cca5"),
                (x"294b39fbd39ce739ce73bdd084a5339ce739ce734a58c9cca5"),
                (x"294b39b5b9cce739ce739cd299ce739ce739a1084a58c9cca5"),
                (x"294b39b5b9cce739ce739cd299ce739ce739a1084a58c9cca5"),
                (x"294b39b5ac656b59ce739ce739ce739ce68421084a58c9cca5"),
                (x"294b39b5ac656b59ce739ce739ce739ce68421084a58c9cca5"),
                (x"294b39b1894a1084a6739ce739ce739a108421084a58c9cca5"),
                (x"294b39b1894a1084a6739ce739ce739a108421084a58c9cca5"),
                (x"294b39b18842108422739ce739ce739a528421084a7399cca5"),
                (x"294b39b18842108422739ce739ce739a528421084a7399cca5"),
                (x"294b39b18842108422739ce739ce739a528421084a7399cca5"),
                (x"294b39b188421089ce739ce739ce739ce694a1084a58c9cca5"),
                (x"294b39b188421089ce739ce739ce739ce694a1084a58c9cca5"),
                (x"294b39e7294ce739ce739cd8c9ce739ce739eb5a631ad9cca5"),
                (x"294b39e7294ce739ce739cd8c9ce739ce739eb5a631ad9cca5"),
                (x"294b39b1939ce739ce739cf39a52939ce739ce73ce5ad9cca5"),
                (x"294b39b1939ce739ce739cf39a52939ce739ce73ce5ad9cca5"),
                (x"294b39ce739ce739cd296318c4a52844e739ce739cd8c9cca5"),
                (x"294b39ce739ce739cd296318c4a52844e739ce739cd8c9cca5"),
                (x"294b39ce739ce739cd296318c4a52844e739ce739cd8c9cca5"),
                (x"294b39ce739ce73ce50842108421094b1939ce739ce739cca5"),
                (x"294b39ce739ce73ce50842108421094b1939ce739ce739cca5"),
                (x"294b39ce739b18c6b58c6318c6318c635ad6ce739ce739cca5"),
                (x"294b39ce739b18c6b58c6318c6318c635ad6ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294b39ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 1719 := 0;
    signal out_color_reg : std_logic_vector(0 to 199) := (others => '0');
begin
    process(in_sprite_id, in_sprite_row, in_sprite_col, in_sprite_state, in_sprite_direction)
    begin
        real_row <= 0;
        case in_sprite_id is
            when 0 => real_row <= in_sprite_row;
            when 1 => real_row <= 40 + in_sprite_row;
            when 2 => real_row <= 80 + in_sprite_row;
            when 3 => real_row <= 120 + in_sprite_row;
            when 4 =>
                case in_sprite_state is
                    when 0 => real_row <= 160 + in_sprite_row;
                    when 1 => real_row <= 200 + in_sprite_row;
                    when others => null;
                end case;
            when 5 =>
                case in_sprite_state is
                    when 0 => real_row <= 240 + in_sprite_row;
                    when 1 => real_row <= 280 + in_sprite_row;
                    when 2 => real_row <= 320 + in_sprite_row;
                    when 3 => real_row <= 360 + in_sprite_row;
                    when others => null;
                end case;
            when 6 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 400 + in_sprite_row;
                            when D_RIGHT => real_row <= 440 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 480 + in_sprite_row;
                            when D_RIGHT => real_row <= 520 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 560 + in_sprite_row;
                            when D_RIGHT => real_row <= 600 + in_sprite_row;
                            when others => null;
                        end case;
                    when 3 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 640 + in_sprite_row;
                            when D_RIGHT => real_row <= 680 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 7 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 720 + in_sprite_row;
                            when D_RIGHT => real_row <= 760 + in_sprite_row;
                            when D_DOWN => real_row <= 800 + in_sprite_row;
                            when D_LEFT => real_row <= 840 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 880 + in_sprite_row;
                            when D_RIGHT => real_row <= 920 + in_sprite_row;
                            when D_DOWN => real_row <= 960 + in_sprite_row;
                            when D_LEFT => real_row <= 1000 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1040 + in_sprite_row;
                            when D_RIGHT => real_row <= 1080 + in_sprite_row;
                            when D_DOWN => real_row <= 1120 + in_sprite_row;
                            when D_LEFT => real_row <= 1160 + in_sprite_row;
                            when others => null;
                        end case;
                    when 3 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1200 + in_sprite_row;
                            when D_RIGHT => real_row <= 1240 + in_sprite_row;
                            when D_DOWN => real_row <= 1280 + in_sprite_row;
                            when D_LEFT => real_row <= 1320 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 8 => real_row <= 1360 + in_sprite_row;
            when 9 => real_row <= 1400 + in_sprite_row;
            when 10 => real_row <= 1440 + in_sprite_row;
            when 11 => real_row <= 1480 + in_sprite_row;
            when 12 => real_row <= 1520 + in_sprite_row;
            when 13 => real_row <= 1560 + in_sprite_row;
            when 14 => real_row <= 1600 + in_sprite_row;
            when 15 => real_row <= 1640 + in_sprite_row;
            when 16 => real_row <= 1680 + in_sprite_row;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= rom(real_row);
        end if;
    end process;
    out_color <= out_color_reg((in_sprite_col * 5) to ((in_sprite_col + 1) * 5) - 1);
end behavioral;
