library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

entity graphic_controller is
    port(
        CLK, RST : in std_logic
        
        
        data_block : in 
    );
end graphic_controller;

architecture behaviorial of graphic_controller is
begin

end architecture;