library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.PROJECT_PARAMS_PKG.all;
use work.PROJECT_TYPES_PKG.all;
use work.PROJECT_DIRECTION_PKG.all;

entity ressources_sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_id : in block_category_type;
        in_sprite_state : in state_type;
        in_sprite_direction : in direction_type;

        in_sprite_row : in integer range 0 to 39;
        in_sprite_col : in integer range 0 to 39;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end ressources_sprite_rom;

architecture behavioral of ressources_sprite_rom is
    subtype word_t is std_logic_vector(0 to 199);
    type memory_t is array(0 to 1679) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- 0_empty
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 1_unbreakable
                (x"ef5ef784210842108421084210842108421084210842318def"),
                (x"ef5ef784210842108421084210842108421084210842318def"),
                (x"ef5ef790810842108421084210842108421084210908318def"),
                (x"ef5ef790810842108421084210842108421084210908318def"),
                (x"ef5ef790810842108421084210842108421084210908318def"),
                (x"ef5ef784210848421084210842108421084210210842318def"),
                (x"ef5ef784210848421084210842108421084210210842318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784242108421084210842108421084210842042318def"),
                (x"ef5ef784210848421084210842108421084210210842318def"),
                (x"ef5ef784210848421084210842108421084210210842318def"),
                (x"ef5ef784210848421084210842108421084210210842318def"),
                (x"ef5ef790810842108421084210842108421084210908318def"),
                (x"ef5ef790810842108421084210842108421084210908318def"),
                (x"ef5ef78c6318c6318c6318c6318c6318c6318c6318c6318def"),
                (x"ef5ef78c6318c6318c6318c6318c6318c6318c6318c6318def"),
                (x"ef5ef78c6318c6318c6318c6318c6318c6318c6318c6318def"),
                (x"ef7def3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef"),
                (x"ef7def3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef"),
                (x"ef7def3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef"),
                (x"ef7bdefbdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde"),
                (x"ef7bdefbdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bde"),
                (x"ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7de"),
                (x"ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7de"),
                (x"ef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7de"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce739c"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce739c"),

                -- 2_unbreakable
                (x"e73bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e73bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e71ef790842108421084210842108421084210842108318fbd"),
                (x"e71ef790842108421084210842108421084210842108318fbd"),
                (x"e71ef790842108421084210842108421084210842108318fbd"),
                (x"e73def0c6108421084210842108421084210842108c6f7bfbd"),
                (x"e73def0c6108421084210842108421084210842108c6f7bfbd"),
                (x"e73def3de1085ef7bdef7bdef7bdef7bdef7bc2108c6f7bfbd"),
                (x"e73def3de1085ef7bdef7bdef7bdef7bdef7bc2108c6f7bfbd"),
                (x"e73def3de1085ef7bdef7bdef7bdef7bdef7bc2108c6f7bfbd"),
                (x"e73def3de108463190842106318c842108f7bc2108c6f7bfbd"),
                (x"e73def3de108463190842106318c842108f7bc2108c6f7bfbd"),
                (x"e73def3de108463190842106318c842108f7bc2108c6f7bfbd"),
                (x"e73def3de1084631bde42106318def7908f7bc2108c6f7bfbd"),
                (x"e73def3de1084631bde42106318def7908f7bc2108c6f7bfbd"),
                (x"e73def3de10846318c6318c6318c6318c6f7bc2108c6f7bfbd"),
                (x"e73def3de10846318c6318c6318c6318c6f7bc2108c6f7bfbd"),
                (x"e73def3de10846318c6318c6318c6318c6f7bc2108c6f7bfbd"),
                (x"e73def3de108463190842106318c842108f7bc2108c6f7bfbd"),
                (x"e73def3de108463190842106318c842108f7bc2108c6f7bfbd"),
                (x"e73def3de1084631bde42106318def7908f7bc2108c6f7bfbd"),
                (x"e73def3de1084631bde42106318def7908f7bc2108c6f7bfbd"),
                (x"e73def3de10846318c6318c6318c6318c6f7bc2108c6f7bfbd"),
                (x"e73def3de10846318c6318c6318c6318c6f7bc2108c6f7bfbd"),
                (x"e73def3de10846318c6318c6318c6318c6f7bc2108c6f7bfbd"),
                (x"e73def3de108421084210842108421084210842108c6f7bfbd"),
                (x"e73def3de108421084210842108421084210842108c6f7bfbd"),
                (x"e73def3de318c6318c6318c6318c6318c6318c6318c6f7bfbd"),
                (x"e73def3de318c6318c6318c6318c6318c6318c6318c6f7bfbd"),
                (x"e73def3de318c6318c6318c6318c6318c6318c6318c6f7bfbd"),
                (x"e73def3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bfbd"),
                (x"e73def3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bfbd"),
                (x"e73def3def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bfbd"),
                (x"e73def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bcf7bfbd"),
                (x"e73def7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bcf7bfbd"),
                (x"e73bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e73bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e73bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bdef7bd"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce73bd"),
                (x"e739ce739ce739ce739ce739ce739ce739ce739ce739ce73bd"),

                -- 3_breakable
                (x"318842108421084210842108421084218c739c6318c6318c63"),
                (x"318842108421084210842108421084218c739c6318c6318c63"),
                (x"39c84210842108421084210842108421ce739c6318c6318c63"),
                (x"39c84210842108421084210842108421ce739c6318c6318c63"),
                (x"39c84210842108421084210842108421ce739c6318c6318c63"),
                (x"39c84210842108421084210842108421ce739c6318c6318c63"),
                (x"39c84210842108421084210842108421ce739c6318c6318c63"),
                (x"39c842108421084210842108421084218c739c6318c6318c63"),
                (x"39c842108421084210842108421084218c739c6318c6318c63"),
                (x"39c842108421084210842108421084218c739c6318c6318c63"),
                (x"39ca5294a5294a5294a5294a5294a5298c739ce739ce739ce7"),
                (x"39ca5294a5294a5294a5294a5294a5298c739ce739ce739ce7"),
                (x"39ca5294a5294a5294a5294a5294a5298c739ce739ce739ce7"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"294a5294a6318a52908421084210842108421084218c318ca5"),
                (x"294a5294a6318a52908421084210842108421084218c318ca5"),
                (x"294a5294a6318a52908421084210842108421084218c318ca5"),
                (x"294a5294a6318a5290842108421084210842108421ce318ca5"),
                (x"294a5294a6318a5290842108421084210842108421ce318ca5"),
                (x"18c6318c6739ca5290842108421084210842108421ce318c63"),
                (x"18c6318c6739ca5290842108421084210842108421ce318c63"),
                (x"18c6318c66318a5294a5294a5294a5294a5294a529ce318c63"),
                (x"18c6318c66318a5294a5294a5294a5294a5294a529ce318c63"),
                (x"18c6318c66318a5294a5294a5294a5294a5294a529ce318c63"),
                (x"39cc6318c6318c631ce6318c6318c6318c6318c631ce739ce7"),
                (x"39cc6318c6318c631ce6318c6318c6318c6318c631ce739ce7"),
                (x"2108421084210842108739c6318c6318c6318cc63108421084"),
                (x"2108421084210842108739c6318c6318c6318cc63108421084"),
                (x"2108421084210842108739c6318c6318c6318cc63108421084"),
                (x"2108421084210842108739c6318c6318c6318cc63108421084"),
                (x"2108421084210842108739c6318c6318c6318cc63108421084"),
                (x"2108421084210842108739c6318c6318c6318cc63108421084"),
                (x"294a5294a5294a5294a739c6318c6318c6318cc6314a5294a5"),
                (x"294a5294a5294a5294a739c6318c6318c6318cc6314a5294a5"),
                (x"39ce739ce739ce739ce739ce739ce739ce739cc631ce739ce7"),
                (x"39ce739ce739ce739ce739ce739ce739ce739cc631ce739ce7"),
                (x"39ce739ce739ce739ce739ce739ce739ce739cc631ce739ce7"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),
                (x"318c6318c6318c6318c6318c6318c6318c6318c6318c6318c6"),

                -- 4_bomb_0
                (x"fffffffffffffffffffffffffffffffffffffffffa11ffffff"),
                (x"fffffffffffffffffffffffffffffffffffffffffa11ffffff"),
                (x"fffffffffffffffffc00000000000000000fffe004e68423ff"),
                (x"fffffffffffffffffc00000000000000000fffe004e68423ff"),
                (x"fffffffffffffffffc00000000000000000fffe004e68423ff"),
                (x"fffffffffff80000039ce739ce739ce73ff0001ff801ffffff"),
                (x"fffffffffff80000039ce739ce739ce73ff0001ff801ffffff"),
                (x"ffffffffe0018c631821318dce739c08400fffe00001ffffff"),
                (x"ffffffffe0018c631821318dce739c08400fffe00001ffffff"),
                (x"ffffff8006346318c631318c63739c084000001ce7380003ff"),
                (x"ffffff8006346318c631318c63739c084000001ce7380003ff"),
                (x"ffffff8006346318c631318c63739c084000001ce7380003ff"),
                (x"ffffff8011884210856b8c6263739cfffffe739ce7380003ff"),
                (x"ffffff8011884210856b8c6263739cfffffe739ce7380003ff"),
                (x"ffc00018d1884210856b8c626318c6e739ce739ce739ce7000"),
                (x"ffc00018d1884210856b8c626318c6e739ce739ce739ce7000"),
                (x"ffc00018d18ad6b5ad6b8c626318c6e739ce739ce739ce7000"),
                (x"ffc00018d18ad6b5ad6b8c626318c6e739ce739ce739ce7000"),
                (x"ffc00018d18ad6b5ad6b8c626318c6e739ce739ce739ce7000"),
                (x"ffc00018d18c6318c6318c626318c6e739ce739ce739ce7000"),
                (x"ffc00018d18c6318c6318c626318c6e739ce739ce739ce7000"),
                (x"ffc00018c6346318c631318c6318c6e739ce739ce739ce7000"),
                (x"ffc00018c6346318c631318c6318c6e739ce739ce739ce7000"),
                (x"ffc00018c6346318c631318c6318c6e739ce739ce739ce7000"),
                (x"ffc0007386318c6318c6318c63739ce739ce739ce739ce7000"),
                (x"ffc0007386318c6318c6318c63739ce739ce739ce739ce7000"),
                (x"ffc000739ce18c6318c6e739ce739ce739ce739ce739ce7000"),
                (x"ffc000739ce18c6318c6e739ce739ce739ce739ce739ce7000"),
                (x"ffffff801ce739ce739ce739ce739ce739ce739ce7380003ff"),
                (x"ffffff801ce739ce739ce739ce739ce739ce739ce7380003ff"),
                (x"ffffff801ce739ce739ce739ce739ce739ce739ce7380003ff"),
                (x"ffffff801ce739ce739ce739ce739ce739ce739ce7380003ff"),
                (x"ffffff801ce739ce739ce739ce739ce739ce739ce7380003ff"),
                (x"ffffffffe00739ce739ce739ce739ce739ce739ce001ffffff"),
                (x"ffffffffe00739ce739ce739ce739ce739ce739ce001ffffff"),
                (x"fffffffffff80000039ce739ce739ce739c0000007ffffffff"),
                (x"fffffffffff80000039ce739ce739ce739c0000007ffffffff"),
                (x"fffffffffff80000039ce739ce739ce739c0000007ffffffff"),
                (x"fffffffffffffffffc00000000000000000fffffffffffffff"),
                (x"fffffffffffffffffc00000000000000000fffffffffffffff"),

                -- 5_explosion_0
                (x"ffffffb339cdb494a538b4e694a6739da79ce739ce7bffffff"),
                (x"ffffffb339ce67ac63189dada4a75ad4ed9ce739ce73ffffff"),
                (x"ffffffe739ce7369ce76b4e694e318c4ed39cf39ce73ffffff"),
                (x"ffffffe739ce7369ce76b4e694e318c4ed39cf39ce73ffffff"),
                (x"fffff66739ce676b5ad3d25294a529d5ad6b6739ce739fffff"),
                (x"f7bde66739cced6b5ada4eb5a4eb5ad4e79ce739ce73963199"),
                (x"7398cce739cced6b5ada4e3094e35a9db39cda73ce739cce6c"),
                (x"7398cce739cced6b5ada4e3094e35a9db39cda73ce739cce6c"),
                (x"eb3399e739ccf33ce678d6b494a673b5a79cdad9ce7399ce6c"),
                (x"ce7399db399cf39ce678d4e7a4a75ad4e739e673ce733b6739"),
                (x"ce739ce673b5ad3ce678c6b584a7184ead6b4e769ce79ce733"),
                (x"ce739cdad6b5a739cf494a5294a5294ead39dad6b5ad39ce76"),
                (x"d6a739dad6b5b589cf5ac25294a5294a7139dad6b5ad6b5ad6"),
                (x"d6a739dad6b5b589cf5ac25294a5294a7139dad6b5ad6b5ad6"),
                (x"4e273b5ad6b4f569cd29d6b49c25294a7539dad6b5a739dad6"),
                (x"4ea73b4ed6b4f56b5b49c21094a5294e2739da769cf18c6b4c"),
                (x"4ea739ce73b5b1ab5a784a1084a5294e27ad6b569cf094a53e"),
                (x"4ead6b5a739cf18d6b5a4a1094a5294e12842709d6b494a53a"),
                (x"4ead6b5a739cf18d6b5a4a1094a5294e12842709d6b494a53a"),
                (x"4a673b5a734a7184a5384a5384a129c250842529d6b49c2538"),
                (x"c612942273c25294a529c63094a1294e3494a53ad693ac2529"),
                (x"4a529425084e1284a749c2528425294ce7ad6a73d6b13d6b49"),
                (x"4a529c6929d61299ce69c252842129427539ce769ce734e309"),
                (x"4a529c6929d61299ce69c252842129427539ce769ce734e309"),
                (x"c275a9dad69a529d6a694a529425294a538c4f13b5ad39a53a"),
                (x"4a75ab5ad69ce7ad6b584a5294e129c25294ea76b5ad9cce78"),
                (x"d4ed6b5ad6b5ad6b5a694a5294a5294a75ad4ed6b5a79b4e7a"),
                (x"9dad6cced6b5ad6b5adad63094a529d4ed6b5ad69cf339ce73"),
                (x"9dad6cced6b5ad6b5adad63094a529d4ed6b5ad69cf339ce73"),
                (x"ce6d69e673b4ed69ced69a538d69299dad6b4ed3ce7369ce76"),
                (x"66739ce739ce739ce733c2538b5a739e676b5a79ce7399ce7e"),
                (x"77739ce739ce739ce7334e31a9ce73d67339e739ce739ce72c"),
                (x"f7739ce739ce673ce73a4a538d6b5ac4ed6b6739ce739ce739"),
                (x"f7739ce739ce673ce73a4a538d6b5ac4ed6b6739ce739ce739"),
                (x"ce73966739ce736b5ad6d25294a529d5ad39e739ce739cb18c"),
                (x"fffff66739ce736b5ad69a5294a75a9dad6b6739ce739fffff"),
                (x"ffffffb339ce736b5ad69ce78422739ce79ce739ce73ffffff"),
                (x"fffffffb39ce736b5ad6b5ad3c275a9cf39ce739ce73ffffff"),
                (x"fffffffb39ce736b5ad6b5ad3c275a9cf39ce739ce73ffffff"),
                (x"ffffff318cce6799cf539dada4250842679ce739ce733fffff"),

                -- 5_explosion_1
                (x"ce7bdf6739ce929c61294a528421084275ad6933b5ad3cfbde"),
                (x"ce58cee6d69a5294a709421084212942538c27539ced3cb199"),
                (x"9dad69ce73d2718c630942108421084a138c6a739ced6ce72c"),
                (x"9dad69ce73d2718c630942108421084a138c6a739ced6ce72c"),
                (x"b5ad6b5a73d61294a52942108421084a53ad6b139ced3ce739"),
                (x"b5ad6b4e739e9294a52842108421084a71ad27139ced69ce73"),
                (x"b5ad6b6b5ad2529c61294a108421084271ad27139ced6b5ad3"),
                (x"b5ad6b6b5ad2529c61294a108421084271ad27139ced6b5ad3"),
                (x"9dad6b4d294a5294a70942108421294a5294a5299ced3b4e73"),
                (x"4ced69db5a4a5294a70942108427184a5294a529d6b49d6b53"),
                (x"4ead6d6b184a718c630942108427184a718c61294a5294eb53"),
                (x"c635ac25294e1294a52842108425294a5294a70942138c2538"),
                (x"4a5294a5294a5294210842108421084210842309421284e309"),
                (x"4a5294a5294a5294210842108421084210842309421284e309"),
                (x"4a529c6129425294210842108421084210842529421084e308"),
                (x"4a1084a5294a1094a5084210842108421084610842109d2523"),
                (x"4a108421084a50942108421084210842108425284210842108"),
                (x"421084210842108421084210842108421094a5084210842108"),
                (x"421084210842108421084210842108421094a5084210842108"),
                (x"42108421084210842108421084210842108421084210842108"),
                (x"421294a5084212842108421084210842108421084210842108"),
                (x"421294a108425384a50842108421294a108421084210842109"),
                (x"463184a1084a5384a50842108421084a1294a5294210842108"),
                (x"463184a1084a5384a50842108421084a1294a5294210842108"),
                (x"4a5294a529421294a5084210842108425294a7184a5384a529"),
                (x"4a5294a5294a1094a5084210842108421294a109c6129c6318"),
                (x"4a529c25294a1184a528421084210842138c2509c61294a529"),
                (x"d61294a718c2538c6309421084210842128461294a5294a529"),
                (x"d61294a718c2538c6309421084210842128461294a5294a529"),
                (x"d69294e1294e3094a529421084210842128427094a529c4e69"),
                (x"4a7184eb184a5294a529421084210842108425294a5294ce78"),
                (x"d6a734e273c2529c63094a5284210842528427184a71a9dad3"),
                (x"9cf5a4e2d6d25384a5384a528421084a5094e3139cf539ce76"),
                (x"9cf5a4e2d6d25384a5384a528421084a5094e3139cf539ce76"),
                (x"b4e739ced69a53a4a5384a108421084a1094a713b5ad6b5ad6"),
                (x"9e6d6b5ad69e313b5b094e3094210842718c6a73b5ad6b4e73"),
                (x"ce6d69dad6b6a739cf494e309421294a5094e313b5a79ce739"),
                (x"ce739cced69ceda4a7094a52842129421094e13ab5b39ce72c"),
                (x"ce739cced69ceda4a7094a52842129421094e13ab5b39ce72c"),
                (x"ce739ce6d6b5b094a7094210842108421094e13ab5b39cf7ae"),

                -- 5_explosion_2
                (x"fe58cce6d69e1284210842108ded0842138c6b1ab599e67bde"),
                (x"fe58cce6d6d21084210842108b8508421294a673b5b2cee72c"),
                (x"cb18cce6739a5294210842108b850842138c2676b5a79ce739"),
                (x"cb18cce6739a5294210842108b850842138c2676b5a79ce739"),
                (x"63339ce718d69294210842108b877b421094e313b5ad99e739"),
                (x"9e739ce718d69284210842108ddef7ba1094a53a9ce76b5ad3"),
                (x"b4f39ceb5a9e9284210845ef7ba1084210842109d6ad69dacc"),
                (x"b4f39ceb5a9e9284210845ef7ba1084210842109d6ad69dacc"),
                (x"b5ad69ea739e92842108b84210ed08425294a1189cf5ac6b4c"),
                (x"9cf5ad6ad6d250842108b8421b86f7421084253ad69284a538"),
                (x"4a50846273c250842108b843746ef742108427494a529c2528"),
                (x"4a108427184210842108def68422f74210846b58c6138c6308"),
                (x"4210842129421084210842117ddef742108461294a5294a529"),
                (x"4210842129421084210842117ddef742108461294a5294a529"),
                (x"4212942108421084210840421ba37b42108425084210842108"),
                (x"421084a508421084210846f61beef7da1094a108421084e308"),
                (x"42108422f7da10842108421080def7da1084237742108c4e68"),
                (x"4210846c21da1084210846f770877b421084237bdef7b42108"),
                (x"4210846c21da1084210846f770877b421084237bdef7b42108"),
                (x"4210846f7bbdd0842108bdee1086f74210842117bdef742108"),
                (x"4210842108bdee84211bba11708421da10842117bdc3742108"),
                (x"42108421084210842108ddefbb86f70a10842108deefb42108"),
                (x"42108421084210842101ba11bbdd084210842108bdefb42108"),
                (x"42108421084210842101ba11bbdd084210842108bdefb42108"),
                (x"4252942108421084a76142117ddd084210842108421084a108"),
                (x"4275a4a108421294a777def7b4237b4210842108421084a523"),
                (x"4a7184a1084213a4a51b0dee8ddd084210842108421094a11e"),
                (x"427184a529c250942108ddef7b877b4210842108421094e31e"),
                (x"427184a529c250942108ddef7b877b4210842108421094e31e"),
                (x"421294a5299e90842108d84210def742108421294a5084631e"),
                (x"9a5084635ad252842108d84210a1084210842318d6b484b18c"),
                (x"b690844e73d21294210845efbda1084210842709d6b5ac672c"),
                (x"b69084dad6d213a4a5084211b421084213ad4f5ad6b53b6739"),
                (x"b69084dad6d213a4a5084211b421084213ad4f5ad6b53b6739"),
                (x"cdb5a9da739a509c612845ee10ed084211ad4e73d6b53b6739"),
                (x"9dad69dad69cd094a51bb8421ba1084a118c4e73c6279b673d"),
                (x"b5ad6b5ad69cf4942361084210a1084a5094a753d6a79ce73e"),
                (x"fcf39b5ad6b4f49422e10843b4210842718c27569ced96319e"),
                (x"fcf39b5ad6b4f49422e10843b4210842718c27569ced96319e"),
                (x"ffd8cce739b6928422e108437bed0842138c2756b5b2c77fff"),

                -- 5_explosion_3
                (x"fffdef318cb250842361084210def7da1294a7569cf2c77fff"),
                (x"fcf39ce7399a5084211bbdee1084210a1084213ad6a7364e73"),
                (x"b4f39cce734a5084210842101086f746d18c2109d6b5ab5ad9"),
                (x"b4f39cce734a5084210842101086f746d18c2109d6b5ab5ad9"),
                (x"b5b39cce734a1084210845ee1bed0845c294a53ad69299ce73"),
                (x"9dad69e9294a1084211bbdee1bdd0845c37ba318c61294a53a"),
                (x"9da73d25294a508422e108421086f7bdee8423094a52842109"),
                (x"9da73d25294a508422e108421086f7bdee8423094a52842109"),
                (x"b4e73d252942528dec21084210842108508421384a5084a529"),
                (x"d69294a5084211b0842108421084210851bda1384a5294e318"),
                (x"4e9294a50842377deef708421084210def7ba138c61294a103"),
                (x"9e9084277b42117ded1708421084210dc210a138421084210e"),
                (x"4a1084210842117ded170842108421bdee10a1094211bbeb59"),
                (x"4a1084210842117ded170842108421bdee10a1094211bbeb59"),
                (x"4a77bba37bddf68dec2108421086f7420210eef7421010def8"),
                (x"4a37b4237bb8437bdc210842108421420210eee1bdef70dee1"),
                (x"46ef7422f70dc210842108421086f746f610df6108768ddee1"),
                (x"45c2108421084210842108421084210842108501086fb46f61"),
                (x"45c2108421084210842108421084210842108501086fb46f61"),
                (x"086f7084210842108421084210842108421087610843746f63"),
                (x"b86f7b842108421084210842108421084210842108421bdeec"),
                (x"46c21bdc210842108421084210842108421084210842108423"),
                (x"4237bb84210dee10842108421084210842108421086e108421"),
                (x"4237bb84210dee10842108421084210842108421086e108421"),
                (x"422f7bdf7bbdd010842108421084210842108437def7bb8421"),
                (x"da108422f70dee1084210842108421086f7beef7bdd0846f77"),
                (x"42108422f7ba2f708421ddee10842108508422f7ded0842108"),
                (x"4210842108aa777bdefb08421084210df77ba2f74210842108"),
                (x"4210842108aa777bdefb08421084210df77ba2f74210842108"),
                (x"4a1084a10842508421170842108421ba2f7ba108421084253e"),
                (x"c6129425294a1084237708437da2f70843bda108421094a109"),
                (x"4a5294ea73c2508bdef7bdef7da2f708437ba10842129c2108"),
                (x"4a5294ce73c2508bdd170ef68422f70dee842528421294ce7a"),
                (x"4a5294ce73c2508bdd170ef68422f70dee842528421294ce7a"),
                (x"c6318d5a734a1084211708437bdef70dd0846b094a5389ce73"),
                (x"cb273d275ad210842117084210def70dd0842509d6b139e739"),
                (x"f7a734a5294a52942361084210dc21bdd08421094a53ace73d"),
                (x"ff7399a52942528bdc210842108421bdd08421384a753ce73f"),
                (x"ff7399a52942528bdc210842108421bdd08421384a753ce73f"),
                (x"fff399a1084251708421084210842108768421299cf39cffff"),

                -- 6_explosion_0_0
                (x"fffffffffff33369cd29c25294a35a9db36b4f39ce7dffffff"),
                (x"ffffffff39ce7369cf094a5294a7189db339cf39633dffffff"),
                (x"ffffffb339cced6b5a7a9eb584a75ab5a76b4f39633fffffff"),
                (x"ffffffb339cced6b5a7a9eb584a75ab5a76b4f39633fffffff"),
                (x"ffffffb339cced39ced6b5ad8d62739da79cced9633fffffff"),
                (x"ffffffb339ce6d3d6b5ad5ac94ce739db39ce7396319ffffff"),
                (x"ffffffb98c9dad69ce73c6b484ce73b5a79ce7396319ffffff"),
                (x"ffffffb98c9dad69ce73c6b484ce73b5a79ce7396319ffffff"),
                (x"ffffffb98c9da76b5ad6d210842673b5b39ce739ce7dffffff"),
                (x"ffffffb98cb6736b5ad34a1084ead69cf339cf39631dffffff"),
                (x"fffffffd8cce676b5ada4a529c4ed69cf36b4f3ef7bfffffff"),
                (x"ffffffff399dad6b5a739a5294ced69dad39e72cf7bfffffff"),
                (x"ffffffdb39ce6d69cd38d630946a739dad39b339633dffffff"),
                (x"ffffffdb39ce6d69cd38d630946a739dad39b339633dffffff"),
                (x"ffffffe739ce676d6929d6b5a4a7189e6739e739ce73ffffff"),
                (x"ffffffe739b5a739cd384e31a4a529d5b39cdad69ce7ffffff"),
                (x"ffffffe739ce6d69ce739eb494a7189da79cdad6ce73ffffff"),
                (x"fffffffb39ce676b5a73d63094a5299dad9ccf39ce73ffffff"),
                (x"fffffffb39ce676b5a73d63094a5299dad9ccf39ce73ffffff"),
                (x"ffffffb339ce736b5ad6c25294a5294da79ce739ce73ffffff"),
                (x"ffffffff39ce7339ce7ac2538c612944ed9ce739ce73ffffff"),
                (x"ffffffff39ce739ce7294a5294e1084cf39ce72cce59ffffff"),
                (x"ffffffb339ce739ce6d3d63094a5294ea79ce72c633fffffff"),
                (x"ffffffb339ce739ce6d3d63094a5294ea79ce72c633fffffff"),
                (x"fffffff98cce6769cf53b63094a7184ead39e72c633fffffff"),
                (x"fffffff98cce6d69cf53b6309c61299da739cf39ce73ffffff"),
                (x"fffffffb39cced69cf53b631a9eb5ab5ad9ccf39ce59ffffff"),
                (x"ffffffb339cced6b5a739a53a9ead6b5ad39e739633dffffff"),
                (x"ffffffb339cced6b5a739a53a9ead6b5ad39e739633dffffff"),
                (x"ffffffb3bd66676b5a76d2109d4e73b5ad9ce739631dffffff"),
                (x"fffffffd8c9e733b5ad3c25294a7189dad9ce72cf7bfffffff"),
                (x"ffffffff399e739b5ad3d6b584a129b5ad9ce73e633fffffff"),
                (x"fffffff7399cf39b5ad6b6b494a1089ced9ce72cce73ffffff"),
                (x"fffffff7399cf39b5ad6b6b494a1089ced9ce72cce73ffffff"),
                (x"ffffffb339cce73b5ad3d253a4a529d5ad39e679633dffffff"),
                (x"ffffffe739cced6b5ad34eb53d27189dad9ce6d3ce7dffffff"),
                (x"ffffffe739ce6d6b5ad6d6b539a7189ce79ce6d6ce59ffffff"),
                (x"ffffffe739ce6769ce769ce73c6273b5ad9ce6d6ce73ffffff"),
                (x"ffffffe739ce6769ce769ce73c6273b5ad9ce6d6ce73ffffff"),
                (x"fffff66739ce6d6d69339eb5a9ce739ce79ce733ce739fffff"),

                -- 6_explosion_0_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"67ffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ce739cb3bdffd8cf7bde67fff67b39ce6dfffdce7398c67fff"),
                (x"ce739ce739cb3b9ce58cce739ce739ce739cb18c63339ce73f"),
                (x"ce739ce739cb3b9ce58cce739ce739ce739cb18c63339ce73f"),
                (x"ce739ce6739cd99ce739ce739ce739b67339e6d39cf39ce73e"),
                (x"ce7399ce73ce7339cf39ce739ce739b6736b6736b5b339e72c"),
                (x"b4ed6b4f39ce676b5ad3ce739cced69ced6b4f33b5ad6b6739"),
                (x"b5ad6b4f39cced6b5ad6ce733b5ad69dad6b5ad6b5a73b5ad6"),
                (x"d4ed6b5ad6b5ad69ce73ce733b5a739ea76b5ad69cf53b4e73"),
                (x"d4ed6b5ad6b5ad69ce73ce733b5a739ea76b5ad69cf53b4e73"),
                (x"4ced6b5ad6b5a73d6b5ab6733b4e734a5339dad69cf569e309"),
                (x"9dad69ced69ced39ce739a53ab4e73c27139ea769cf56d2529"),
                (x"9cf5a4ead6d6353b5ad6d2538c6a734eb539a53ac63569a538"),
                (x"d4f5ad275ad2509c6318c25294e35ac6b094a508d6ad6d2529"),
                (x"d4f5ad275ad2509c6318c25294e35ac6b094a508d6ad6d2529"),
                (x"d4e739e929c253ad69294a5384a529d69294a50842138c2529"),
                (x"9e273d25294a7539cf094a5384a5294a5094e1284a53a4a529"),
                (x"9e1294a5084267ad6b094e3184a5294a7539cf499ce784a528"),
                (x"9cf18c25084e276d69384a1094a7184e276b5ad39ce73d631a"),
                (x"9cf18c25084e276d69384a1094a7184e276b5ad39ce73d631a"),
                (x"9da739ea73b4ed6b5a694a5284ce73d4e739ce76b5a73b4e73"),
                (x"9da73b5a73b5ad6b5adad4e73b5ad6b66d6b4e76b5ad6b5ad6"),
                (x"9da73b5ad6b5ad6b5a769e7369da73cced6b67399cf339e739"),
                (x"ce739ccf39ce733ce673ce739ce739cce739da79ce739b4e76"),
                (x"ce739ccf39ce733ce673ce739ce739cce739da79ce739b4e76"),
                (x"ce739ce739ce7399ce79ce739cced6b6599cce79ce7339ce73"),
                (x"cdad6b4f39ce739ce739ce739ce6d6b6739ce739ce736ce739"),
                (x"9dad69e58cf3339ce72c63199ce6d6b672c67b39ce739ce739"),
                (x"ce739cb3396798cce72c66739ce7399e59ef79996318c63199"),
                (x"ce739cb3396798cce72c66739ce7399e59ef79996318c63199"),
                (x"ce58cf7b39ffdde6333ffb199ce7399e7dfffdde6319fffbde"),
                (x"cfffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 6_explosion_1_0
                (x"fffde666739ced3c61389ce7ad69294a759ce739ce73967fff"),
                (x"fff39cced6b5ad34a529d4e694a5084253ad5a739cf39cffff"),
                (x"fff39ce7399dada4a708421084a10842718c6a76b5b39cffff"),
                (x"fff39ce7399dada4a708421084a10842718c6a76b5b39cffff"),
                (x"ffd8c66739cdad34a5284210942108427139cf539cf39cffff"),
                (x"fffffce739cdad69cd28425294a5294a3139cf539cf39cffff"),
                (x"fffffeb3399dad3d6928421094a508423539eb59ce73967fff"),
                (x"fffffeb3399dad3d6928421094a508423539eb59ce73967fff"),
                (x"fffdef318c9cf494a52942108421084a75ad6356ce72c67fff"),
                (x"ffdce64f399e129c61294a5284275ac27539eb56b5b3d77fff"),
                (x"fffff65ad69a529c612842108427184a75ad6a739cf2cfffff"),
                (x"fffff64ed6b6138c6128421084e1294a5294ea76b5ad9fffff"),
                (x"ffdce666d6b693ac6129421094a5294a5294a756b5ad3cffff"),
                (x"ffdce666d6b693ac6129421094a5294a5294a756b5ad3cffff"),
                (x"fffbdce6739eb53d6929421084a5294a538c4ed69ce73cffff"),
                (x"fff39cda73d4ed6d6908421084a529c613ad4f539cf39cffff"),
                (x"fffdef66d6b4e73d69284210842529d61294a533b5ad9effff"),
                (x"fffdef6739b5a73d6b584a108421084a5294a716b5a7967fff"),
                (x"fffdef6739b5a73d6b584a108421084a5294a716b5a7967fff"),
                (x"fffbd66673cda7ad6b094a108421294a5294a713ce73967fff"),
                (x"ffdce66673b5ad69cf0942108421084e1294eb13b5b39cffff"),
                (x"fffbdce739cce73b5b494a108421084a5294ce73b5ad9cffff"),
                (x"ffd8cce739ccf539cf494a109421294a5294ced69ced9cffff"),
                (x"ffd8cce739ccf539cf494a109421294a5294ced69ced9cffff"),
                (x"fff39cb3399da7ad69384a10842108425294ea739ced3cffff"),
                (x"fffff63273b5a7a4a53842108421084275ad6b1ab5ad3cffff"),
                (x"fffffee6d69ce694a7094a108423184e35ad4f1ab5ad3cffff"),
                (x"fffdef33399e129c6129d2528423184a7539ea79ce739cffff"),
                (x"fffdef33399e129c6129d2528423184a7539ea79ce739cffff"),
                (x"ffd8c6798cb69294a5294a528421294a5294ead9ce739cffff"),
                (x"fffff733399ea7a4a5084210842129c25294ead6ce739fffff"),
                (x"fffff733399a676d6929421094a129c26739ced3ce72cfffff"),
                (x"ffe7373273b27569cd29421094a7184e2d39ead6ce58ef7fff"),
                (x"ffe7373273b27569cd29421094a7184e2d39ead6ce58ef7fff"),
                (x"ffd8c666d69a6769cf4942108421294e358c6276b5b2c67fff"),
                (x"fffbdcda739dad3c63484210842108427094ea799ced9cffff"),
                (x"fff399dad6b4e7a4a5294210842108425294e279ce739cffff"),
                (x"fff399e7399cf494a50942108421084a7094ead6b5a7967fff"),
                (x"fff399e7399cf494a50942108421084a7094ead6b5a7967fff"),
                (x"f3339ce673c61294210842108421294e1294ced6b5ad367fff"),

                -- 6_explosion_1_1
                (x"f7ffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"67ffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ce739eb273ffd9effff9677aeefbdecf5dfffddefffecce73e"),
                (x"ce739eb273ffd9effff9677aeefbdecf5dfffddefffecce73e"),
                (x"cce73cb1ce7399eef599ce72c67bdece58c6319eef72cce72c"),
                (x"ce6d6b658c633ccce58cce739ce739b67339da6c63339cce79"),
                (x"9e6d69da73ce599b5a79ce7339e6d69ced6b5b2cce739cdad3"),
                (x"9e6d69da73ce599b5a79ce7339e6d69ced6b5b2cce739cdad3"),
                (x"c4ed69ced69ced39ced3ce736cdad6d4ed6b4e739cf399dad3"),
                (x"c4e73b25294eb589ced69ce76b5a739eb58c2713b5ad6b5ad3"),
                (x"4ea73b4f5a9cd299ce73d4e769ce73b69294a53ab5ad6b5ad6"),
                (x"4a75a9dad6b69294a75a9ce76d4e73b4f58c25299ced3d4e73"),
                (x"42529c4e73d25384a53a9dad3d6b5ad6b18c6309d6a694a538"),
                (x"42529c4e73d25384a53a9dad3d6b5ad6b18c6309d6a694a538"),
                (x"42129d69294a129c6129d6b58c6929425294a5294a529c2529"),
                (x"42529425294a1294a7184a5294e10842528421294210842538"),
                (x"42108421084213a4a5094a5284a50842108421284210846b53"),
                (x"42108421084212942108421084210842108421284212844e73"),
                (x"42108421084212942108421084210842108421284212844e73"),
                (x"42108421294a108421084a1084210842128421084a5294253a"),
                (x"42108421294a1084210842108421084a5294a1084a5284a53a"),
                (x"4210842129421084210842108421294a538c25284a5284253a"),
                (x"4a108427184a538c61084a1084a1294a5294e3484212842109"),
                (x"4a108427184a538c61084a1084a1294a5294e3484212842109"),
                (x"4a50842529c61294a5084a5294a75ac25294a7094212842109"),
                (x"c25294e3184a529c61294a5384a718c25294a529421094a529"),
                (x"4e129c6ad69a53ad6b494a5294a5294a5294eb5ad6b18c253a"),
                (x"4a5294e2739a533d6b494a5294a529d61294ea7a9ce73c6b59"),
                (x"4a5294e2739a533d6b494a5294a529d61294ea7a9ce73c6b59"),
                (x"9eb18d635a9eb5a9cf5a9ce7a4a5299cd3ad6b58d6a73d5ad9"),
                (x"b5a739ced6b5ad3c6313b4e78c6129d5b539cf5ad6b5a9ce79"),
                (x"b5b39cdad69db39d6b53b4e739da739dad6b4ed6ce673b4e79"),
                (x"b5b399db39ce739b5ad39dad6cdad69ced6b4ed9ce673b4e79"),
                (x"b5b399db39ce739b5ad39dad6cdad69ced6b4ed9ce673b4e79"),
                (x"b4f39b658cce739b5ad6b5ad9cced6cced6b6739ce739ce739"),
                (x"9e739cb1ce667399ce73ce739ce739cce79cb3acce739ce739"),
                (x"63339cb3defff39ce739ce739633bdce73fffdcc63339ce72c"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 6_explosion_2_0
                (x"fb18ccced69e1284a508def77da1084a7494a753b5ad6cfbdf"),
                (x"fb339cced69ea784a50846f61ba1084a7494a75a9ced69b19f"),
                (x"fe739cced6b4e7a4a50842117b86f742108427539cf56ce73f"),
                (x"fe739cced6b4e7a4a50842117b86f742108427539cf56ce73f"),
                (x"fb18ccdad6b69384210846f77bdc21ba10842109c6356cb19f"),
                (x"ffbbd65ad69e129421084211bb877b42108421094a676639df"),
                (x"ffffff4ed6b69294210842117b85084210842753b5ad6639df"),
                (x"ffffff4ed6b69294210842117b85084210842753b5ad6639df"),
                (x"ffffff6673b5b484210842108d8508421084213ab5ad967fff"),
                (x"fb3deee6d6b5a68421294210845f7bda10846b5ab5ad9f7fff"),
                (x"fa58cce6d6b4e784212845efb4237bba118c4ed3b5accf673f"),
                (x"fa273cdad69e128421284042108421bed0842753d6a6ccce7f"),
                (x"fa339cce739a5284210840421084210dd084213a9ce79ce73f"),
                (x"fa339cce739a5284210840421084210dd084213a9ce79ce73f"),
                (x"fa0636335a9cf49c610845ef7b86f7bed094a113b5a6ccb19f"),
                (x"fa35ad6673d5a7ac6128d84370877b421094a6769cf39cfbdf"),
                (x"fe339b6673b5a694a52845ee1bdd0842128426d6b5ad9cfbdf"),
                (x"fe339ce7399da784210845ef7ded084252844ed3b5ad9639df"),
                (x"fe339ce7399da784210845ef7ded084252844ed3b5ad9639df"),
                (x"fa339ce739cdada4212942117da1084271ad4ed3b5ad9cb19f"),
                (x"fe339ce739ccf484212842108bdd08425294ce7a9ce79ce73f"),
                (x"feb39b5a739e9084a52946f61bdef7da12842349d6a79ce73f"),
                (x"fe18ccda73b59294210842108b8421bed094a1339ce79ce73f"),
                (x"fe18ccda73b59294210842108b8421bed094a1339ce79ce73f"),
                (x"fa7bdce673b4f484210846f77beef7da10842356b5b39ce73f"),
                (x"fbbbdce673b69284210846f61ba10842108426769ce79ce73f"),
                (x"fffff666d6b4d284210846f7b421084210842353ce72cb673f"),
                (x"ffffff7b39b5b4842108421084237bda1094a67ac633d9ffff"),
                (x"ffffff7b39b5b4842108421084237bda1094a67ac633d9ffff"),
                (x"ff98c63273b4e694a52942108b86f742118c4e7a4a66c77fff"),
                (x"ff98cf6673b69294a5284211bbdf7b4211ad4f569cf53677bf"),
                (x"fe739cced69a7084210842108bdef742118c5a739cf53cb19f"),
                (x"fcf399dad69ce694212842108b877b421094ce739ce76b319f"),
                (x"fcf399dad69ce694212842108b877b421094ce739ce76b319f"),
                (x"fced6b5ad69da694a50942108b8508425294a533b5ad6b673f"),
                (x"fe6739da73d5b494a5084211b0df7b4e1294a533ce6799e73f"),
                (x"ffb39ce6734ce73d692842101bdf7b425294a51ace739ce73f"),
                (x"ffb39ce6739ea769cf4945ee1bed084270842109b5a79ce73f"),
                (x"ffb39ce6739ea769cf4945ee1bed084270842109b5a79ce73f"),
                (x"fced6b4ed6b4e769cf0845ee84210842718c25094a539ce73d"),

                -- 6_explosion_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"9fbdecce73cfbdfffdc9c6b5846318421084259ffffcccb18c"),
                (x"b67399db39cb19ffffbd66739ce739d0f339b3dffffacce72c"),
                (x"b67399db39cb19ffffbd66739ce739d0f339b3dffffacce72c"),
                (x"b67399da73cf99e63339cdad9ce6d6d3339ce7bef7999ce739"),
                (x"9e739b5ad69e59ece739b5ad9ce739cb276b67399ced69ce73"),
                (x"b4e739dad6b4e79b5a739ce79ce6739ea76b5ad3b5ad6b5ad6"),
                (x"b4e739dad6b4e79b5a739ce79ce6739ea76b5ad3b5ad6b5ad6"),
                (x"b4d29d4e739dad6b5ad6b4e79cced6d4e739dad6b5a76b4e73"),
                (x"9ea73b5a734ea769cf53b6b53b5ad6b4d38c4ed6d6b1a9eb58"),
                (x"9ce73d4e73c267a4a53a4a11ab4e739e9294ce7a4a5299ce69"),
                (x"b5a734a52942528421084a108d6129d2508461084a538d6308"),
                (x"9cf5a4a50842528421084252842129c610842108421084a529"),
                (x"9cf5a4a50842528421084252842129c610842108421084a529"),
                (x"c6929421294252842108425294a1294a1094a5284210842108"),
                (x"42508425084212842108425284a10842108421284210842108"),
                (x"421084210842108421084210842108da10842108421084211b"),
                (x"bdd084210842108def7b46f6845ef70dc210dd084211b46f7b"),
                (x"bdd084210842108def7b46f6845ef70dc210dd084211b46f7b"),
                (x"40421da10846d08dec3740428bdc21bdc210ed08bdf77b8437"),
                (x"45ef70def7bdee8422f7bdef7deef70dc210a11bbdef7bdefb"),
                (x"46ef7b8421bdc284211b0def746ef7084210a2e1084370a108"),
                (x"4237bda37bbeefb421170dee842108ddc210ef6842361ba108"),
                (x"4237bda37bbeefb421170dee842108ddc210ef6842361ba108"),
                (x"421084a1084211b4211bbef684210845c37bdf684211742529"),
                (x"4a529c25084210842108da1094a50846efbda1084210842529"),
                (x"c61294a508421084210842529c252942108421084210846b5a"),
                (x"c21294a529c6b09421084a109d21084a508461084210842529"),
                (x"c21294a529c6b09421084a109d21084a508461084210842529"),
                (x"4a1294a673b4e6942128421139cd294a1094cf484a5084a529"),
                (x"421084a6739ea73d6a7a4eb53b5ad69a13ad5b49d6908d6b5a"),
                (x"4a75a9ce739db5a9ced69a53a9ced6b4f539cf5a9cd299eb53"),
                (x"4db39cda739cd38ce6769eb53b5ad69da7ad5ad6b59389ce76"),
                (x"4db39cda739cd38ce6769eb53b5ad69da7ad5ad6b59389ce76"),
                (x"4cf399da73d6a79ce6799ce73b5ad6cce739dad6b5a7ad5ad6"),
                (x"ce739cdad69cd9d63339ce739ce739cb32c63339b5ad6b5ad6"),
                (x"ce7399dad6cb1d3b5b39ce739cb339ce739cfbcc63199cce79"),
                (x"ce739ce58c677ffce739ce73963bdef33339e7ff739cccb19e"),
                (x"ce739ce58c677ffce739ce73963bdef33339e7ff739cccb19e"),
                (x"f7ffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 6_explosion_3_0
                (x"b4e73b5ad6b5ad34a50842108421084253ad21084a673cb18c"),
                (x"667399ced69ce7a4a51bb843b4237bda10842108421299e739"),
                (x"ef98c9da734a108423610843b45c21ba108425094a53ace73f"),
                (x"ef98c9da734a108423610843b45c21ba108425094a53ace73f"),
                (x"ffd8cce6734a108422b70def7b8421bed294a518d6b53cffff"),
                (x"fffbdce75a4a50842108bef61084210dd08425189ced3cffff"),
                (x"fff39b675a425294a508b84210dc210876842538b5b39cb19f"),
                (x"fff39b675a425294a508b84210dc210876842538b5b39cb19f"),
                (x"ffd8cb5a73425094a53bb843bbdc21086e8421389ced3cfbce"),
                (x"ffe73b5a734e129421080defb08421bdd08421299ced6cb18c"),
                (x"ffed6b5a734a70942108d8421b8421ba1084211ab5ad6b4e79"),
                (x"65a73d4f5ac25294211bb8421bec21ba368421099ce73ce739"),
                (x"cce73d25294a1084211708421da2f7086e8421084a759ce73f"),
                (x"cce73d25294a1084211708421da2f7086e8421084a759ce73f"),
                (x"ce6d69a52942108421170842108421ba10842109d6ad6b7fff"),
                (x"d66d6d2718421284236108421b86f70ed0842129d6ad6b7fff"),
                (x"ce6d69ea73c25284236108421b8508ded08421389ced6b7fff"),
                (x"b6739b5ad6d21284211b0def7bdef74210842529d6b53b7fff"),
                (x"b6739b5ad6d21284211b0def7bdef74210842529d6b53b7fff"),
                (x"64f39b5a73c2529deefbba10846ef7da10842529d6b539e73d"),
                (x"cced69dad6d21084236842108ddf7b4210842108d6a76cb18c"),
                (x"ce739cced6d21084210845efbbdef742508421099ce7963199"),
                (x"d3339cda73d25084211bb84210ec2142528421099ce73f319f"),
                (x"d3339cda73d25084211bb84210ec2142528421099ce73f319f"),
                (x"fff39cdad64a1084236108421dec21da1094a528d6a739ffff"),
                (x"fff399ce734210842108bdefbddc21ba1084271ac6273cffff"),
                (x"fff5ac25084250842108def7708421ba1294e129c6273cb19f"),
                (x"ffd294a50842108422f7bdee1086f7da1294e3099cf39ce739"),
                (x"ffd294a50842108422f7bdee1086f7da1294e3099cf39ce739"),
                (x"ffe739cf5a42108423610dee1bdf7bda1084253a9ced3ce739"),
                (x"ffed6b5a73c25084236108421da2f7ba10842109b5ad3ce72c"),
                (x"1b2d6b5ad69a508422e1084210877b0ed08421089ced667bde"),
                (x"d76d6b4ed6d250842117084210877b0ed0842109b5a76f7bcc"),
                (x"d76d6b4ed6d250842117084210877b0ed0842109b5a76f7bcc"),
                (x"ce6d69ce73c211bbdee108421086f7ba108421089ce7367fff"),
                (x"ce673b5b184a11b08421ddee1084210dd0842108c6279effff"),
                (x"f7739b4d2942508dec21b843b084210dee8421299ce6c77fff"),
                (x"fb98cccd29d2508422e1bdefb406f74210842138d6a79cffff"),
                (x"fb98cccd29d2508422e1bdefb406f74210842138d6a79cffff"),
                (x"ffd8ceb35a9a508422fb46f7b45ef742108421384a713b7fff"),

                -- 6_explosion_3_1
                (x"fffdece75a1fffffffffd673965b39d672c67ffffffffeb196"),
                (x"fbbbdce7bd67ffffffff667339e739ce676b7fffffffff6733"),
                (x"633399dad6b5a69d6b39ce736ce6d6b5a739da6cce7ac66733"),
                (x"633399dad6b5a69d6b39ce736ce6d6b5a739da6cce7ac66733"),
                (x"ee6d6b4ed6b5a69c6279ce733b5a73d4f5ad5ad6b5b399ce76"),
                (x"64e73b4e73b5a694a676b4e76b5b5a4a5339dad6ce739b4e76"),
                (x"d2529c4ed6b4f48422769dad69da73c253ad4e73d6b539dad6"),
                (x"d2529c4ed6b4f48422769dad69da73c253ad4e73d6b539dad6"),
                (x"9e9084e35a9e10842109d6b5ac6b1842138c2528421294ce76"),
                (x"4a529421294a5084a5084a1084a129421094a7094a52844e76"),
                (x"42108421084210842108421084a5294a1094e1284a50844e76"),
                (x"42108ded084210842108421084a108421094a5294a50846b53"),
                (x"4237b0dd08421084210842108da10842108421094a50842529"),
                (x"4237b0dd08421084210842108da10842108421094a50842529"),
                (x"bdc210dd08bef774211b4211bba37bda1084210942115da108"),
                (x"d8421086f70843742101da108dec210defbda11b421170ef68"),
                (x"45ef7d842108437deee1ba108b842108437bec37bdee10dee8"),
                (x"ddc21b8421086f7deee10dee845c2108421086e10877708428"),
                (x"ddc21b8421086f7deee10dee845c2108421086e10877708428"),
                (x"def7b0842108421bdf610ef6845c21084210877b08437def68"),
                (x"42021084210eee10877b0defb45ef7b8777bdc370843742108"),
                (x"b8421084210a2e1086fbddef7ddc210851bd8437bdc21ba108"),
                (x"bdc210df7bddf77084210defbbdd08b86e108421084210ef68"),
                (x"bdc210df7bddf77084210defbbdd08b86e108421084210ef68"),
                (x"420210dc210df7bbdefb42108da37b0dc37bdee108437bef68"),
                (x"422f7ba37bda108421084a5284237bda028422e1086fb42109"),
                (x"422f742108421094a5084a10842108422fbda117ded0942109"),
                (x"4210842108421094a50942108421084210842108421094211a"),
                (x"4210842108421094a50942108421084210842108421094211a"),
                (x"421084210842138c6129421084a50842108421084a5294a108"),
                (x"4a52942108421384a709421084a5294a108421294a50842108"),
                (x"c612942129427494a7484a5284a7184a5094e938c63184a108"),
                (x"4ea73c4ed69da73c631a9ce7ad6a73d69339da73b5a7a4a109"),
                (x"4ea73c4ed69da73c631a9ce7ad6a73d69339da73b5a7a4a109"),
                (x"c4e739ce73b5ad99ce739ce73d6ad6b5b539dad6ce6da4a533"),
                (x"9e58ccced6b4e799ce739e7369ced6b5b339dad3ce673d2533"),
                (x"b65ceeb3de66739ce733f31999dad6b5b39cdb39ce739cce79"),
                (x"ffffffffdef6739633ff6318ccfffffff39ccd9e633ffce72c"),
                (x"ffffffffdef6739633ff6318ccfffffff39ccd9e633ffce72c"),
                (x"fffffffd8cf3339ffffffe72ceffffffff9ce58effffffe72c"),

                -- 7_explosion_0_0
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffe6672cce739cfffffffffffffffffff"),
                (x"fffffffffffffffffffe6672cce739cfffffffffffffffffff"),
                (x"ffffffffffffffffff39ce739ce739ce7fffffffffffffffff"),
                (x"fffffffffffff39ce739ce739ce739ce739cb3ffffffffffff"),
                (x"fffffffffffe7399cf39ce739ce6739e739cb19fffffffffff"),
                (x"fffffffffffe7399cf39ce739ce6739e739cb19fffffffffff"),
                (x"fffffffffff6739b5b39ce739ce6739da79ce739ffffffffff"),
                (x"ffffffffff66733ce739ce739cdad6b5a79ce739ffffffffff"),
                (x"ffffffffffce673ce679cce79cda739cf39ce739ffffffffff"),
                (x"fffffffd8cce739b5b39cce739e673cce79ce739633fffffff"),
                (x"ffffffb18cce7399ce79cdad6b5ad6cce76b5b39631dffffff"),
                (x"ffffffb18cce7399ce79cdad6b5ad6cce76b5b39631dffffff"),
                (x"ffffffe739ce7399ce76cdad6b5ad6b5ad6b4f39ce7bffffff"),
                (x"ffffffb339ce739ce6769eb53b4e73b5ad6b4f39ce59ffffff"),
                (x"ffffffe739ce6799cf56d2529c2673b5ad39e739ce59ffffff"),
                (x"ffffffe739ce733b5a76d25384a75a9da79ce739ce7fffffff"),
                (x"ffffffe739ce733b5a76d25384a75a9da79ce739ce7fffffff"),
                (x"ffffffe739ce7399ced3c25294e9294ea79ce739ce7fffffff"),
                (x"ffffffff39ce739ce6d3c25294ea73d6a739cf39ce7bffffff"),
                (x"ffffffff39cda79b5ad34a53a9dad6b5a739dad6ce7bffffff"),
                (x"ffffffe7399dad9b5ada4a53a9ea73b4f539da73ce59ffffff"),
                (x"ffffffe7399dad9b5ada4a53a9ea73b4f539da73ce59ffffff"),
                (x"ffffffe7399dad6b5ad3d2533d635a9ced39e739ce59ffffff"),
                (x"ffffffe739cdad6b5adad6b53d4f5a4ced9ce739ce59ffffff"),
                (x"ffffffb339ce6d6b5ad3c4e73d4e739dad39e739ce73ffffff"),
                (x"ffffffffdece736b5ad69ce784a6739ced6b6739ce7fffffff"),
                (x"ffffffffdece736b5ad69ce784a6739ced6b6739ce7fffffff"),
                (x"fffffffdcef33399ced6b63094e2739ced6b6739633fffffff"),
                (x"fffffffbdef7b399ced69a5294e273d4e739da79ef7dffffff"),
                (x"fffffffbdece7339ced3c2529d6b5a9ce739dad9f7bdffffff"),
                (x"fffffff98cce6769ced6d2538d6318d4e739cf396319ffffff"),
                (x"fffffff98cce6769ced6d2538d6318d4e739cf396319ffffff"),
                (x"ffffffb98cce676b5a739eb58d6b5ad6b539ce79ce73ffffff"),
                (x"ffffffb98c666769cf53b6b49d6b18c6b539ce6cf7bbffffff"),
                (x"ffffff7bdece736b5a769e3094ea73d6b1ad4e796319ffffff"),
                (x"ffffffb98cce6739ce769eb49c6b5ad4f5ad4e79ce73ffffff"),
                (x"ffffffb98cce6739ce769eb49c6b5ad4f5ad4e79ce73ffffff"),
                (x"ffffffb98cce72c9ce739eb5ac6b5a9ce739cf3ef7bbffffff"),

                -- 7_explosion_0_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffdefffffffffffffffffffffffffffffffffffffffffffff"),
                (x"73bde73bdef7bff63339cffffce7396659ffffffffffffffff"),
                (x"633de6318cf79dece739ce739ce739ce58c67fffffffffffff"),
                (x"633de6318cf79dece739ce739ce739ce58c67fffffffffffff"),
                (x"ce73966739cfbd9ce7339e739ce739ce739ce59effffffffff"),
                (x"ce739ce739cf999ce6d6b5ad9ce739ce739ce739ce7fffffff"),
                (x"ccf399ce73ce739b5ad6b4e79ce673ce739ccf39ce73ffffff"),
                (x"64ed6b5ad69e736b5ad6ce739ccf39ce739cce79ce73ffffff"),
                (x"9ced69da739ce76b5ad6b5ad99da73cce76b67369cf3ffffff"),
                (x"9ced69da739ce76b5ad6b5ad99da73cce76b67369cf3ffffff"),
                (x"9ce73d4ed6b5ad6b5ad6b5ad6b4f5a9ce79ccf39ce739fffff"),
                (x"9dad69ced69dad69cf53d4e739dad6b5b39ce739ce739f7fff"),
                (x"9ce73b4f5ac4ed3c635a4a538c6b5a9e739ce739ce73967fff"),
                (x"d6b18d69294a7139cf494a5294a529d5ad39cf39ce739cffff"),
                (x"d6b18d69294a7139cf494a5294a529d5ad39cf39ce739cffff"),
                (x"d25294e3184a5389ce73d6b494e1299dad39e739ce73967fff"),
                (x"c6129d6b5ad2529d6b5a9ce694a718b5ad39e739ce739cffff"),
                (x"d6b5ad6b18d63099ce78d5adad25299dad9cdad9ce739cffff"),
                (x"d6a73c6b18d4e739cf5a9dad34ea739dad39ced39cf39cffff"),
                (x"d6a73c6b18d4e739cf5a9dad34ea739dad39ced39cf39cffff"),
                (x"9eb5ac6b5a9ea739cd33b5ada4ced6b5b39cced39cf39cffff"),
                (x"9cf5ad6a739ce73b5a739dadad5ad6b5a739ced6ce739fffff"),
                (x"9eb18d6a739ced6b5ad6d4e739ced6b5a739e673ce73ffffff"),
                (x"9eb5a9ce739ced69cf339ce73ce673b5ad9ce739ce73ffffff"),
                (x"9eb5a9ce739ced69cf339ce73ce673b5ad9ce739ce73ffffff"),
                (x"9ce739ce73b5b39ce739b5ad3ce7399ced9ce7396319ffffff"),
                (x"cce739cf39b4f39ce7399dad9ce739ce739ce739633fffffff"),
                (x"f673966739ce739ce7399dad9ce739ce739ce739ffffffffff"),
                (x"f658cf658cf7599ce739ce739ce739ce58c67fffffffffffff"),
                (x"f658cf658cf7599ce739ce739ce739ce58c67fffffffffffff"),
                (x"ee58cee58cf7bffce58c677bdffd8c675dffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_0_2
                (x"fffffff7def66739ce73d6b58d6a739ce6c66739631dffffff"),
                (x"ffffffe739cce7ad6a7ad6b584ea73b4e739cf39631dffffff"),
                (x"ffffffb18ccce7ac635a9eb494e273b4ed6b6739f7bdefffff"),
                (x"ffffffb18ccce7ac635a9eb494e273b4ed6b6739f7bdefffff"),
                (x"fffffff7de64e73d6b58c6b5a4ead69ea76b4f2c631dffffff"),
                (x"ffffffe739cce73d6b5ad6b5ac6a739ced6b4f39631dffffff"),
                (x"ffffffb18cce6739ce7ac631ac275ab5a76b4f39633dffffff"),
                (x"ffffffb18cce6739ce7ac631ac275ab5a76b4f39633dffffff"),
                (x"fffffffbdecdad39ce73d6b5a4a7189da739e739f7bdffffff"),
                (x"fffffffbbdcced39ce7a9e3094a673b5a79ce7def7bdffffff"),
                (x"fffffffd8cce736b5a739e3094e2d6b5a79ce59e73bfffffff"),
                (x"ffffffff39ce736b5a739a529c4e73b5ad6b6739f7bfffffff"),
                (x"ffffffe739ce733b5ad39ce7a9cf189dad6b5b39ce59ffffff"),
                (x"ffffffe739ce733b5ad39ce7a9cf189dad6b5b39ce59ffffff"),
                (x"ffffffb339ce739b5a69d4e7a9eb5ad5ad6b5ad9ce73ffffff"),
                (x"ffffffb339ce733b5a73d631a9a75a9dad6b5ad3ce73ffffff"),
                (x"ffffffb3399ced3d6a769eb53d2529d5ad9cdad3ce73ffffff"),
                (x"fffffff739b5ad39ced6b5ad3d25299dad9cced9ce7fffffff"),
                (x"fffffff739b5ad39ced6b5ad3d25299dad9cced9ce7fffffff"),
                (x"fffffff739ce6739cf5a9eb494a7189db39ce739ce7fffffff"),
                (x"ffffffff39ce7399cf494eb494a7189da79ce739ce73ffffff"),
                (x"ffffffff39ce7399ced3d2529c275ab4ed39e739ce73ffffff"),
                (x"ffffffb339ce733b5ad69a5384a75ab6a79ccf39ce73ffffff"),
                (x"ffffffb339ce733b5ad69a5384a75ab6a79ccf39ce73ffffff"),
                (x"ffffffb339ce676b5ad69ce769ea73b4f39ce739ce59ffffff"),
                (x"fffffff739ce676b5ad6b5ad6b5b39b4e79ce739ce73ffffff"),
                (x"ffffffb98cce6d69ce79b5ad6b5b39cce79ce7396319ffffff"),
                (x"fffffffd8cce7399ce799e7339cf39ce6d9ce739633fffffff"),
                (x"fffffffd8cce7399ce799e7339cf39ce6d9ce739633fffffff"),
                (x"ffffffffffce739ce6739dad9ccf39ccf339cf39ffffffffff"),
                (x"ffffffffffce7399ced6b5ad9ce739ce7339e72cffffffffff"),
                (x"ffffffffffce7399ced39e739ce739ce6d9ce73effffffffff"),
                (x"fffffffffffb199ce7339e739ce739ce679ce73fffffffffff"),
                (x"fffffffffffb199ce7339e739ce739ce679ce73fffffffffff"),
                (x"ffffffffffffd99ce739ce739ce739ce739ce7ffffffffffff"),
                (x"ffffffffffffffffff39ce739ce739ce7fffffffffffffffff"),
                (x"fffffffffffffffffff9ce7396658cf7ffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_0_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff73bac67fffef58c6333ffffde6333d6673d"),
                (x"fffffffffffffec63339ce739ce739ce739cb3be6333e6673e"),
                (x"fffffffffffffec63339ce739ce739ce739cb3be6333e6673e"),
                (x"ffffffffffce739ce739ce739cda73ce739ce739ce72cce73e"),
                (x"fffffffd8cce739ce739ce739cda73ce739ce676ce6739ce79"),
                (x"ffffffb18cce739b5a73ce7399dad6ce739ce6d69ce739ce73"),
                (x"ffffffe739ce739b5ad69e7399ce739e676b5a739ce73d6b53"),
                (x"ffffffe7399cf339ced6b4e739cf5ab5ad6b5a739cf5ac6b53"),
                (x"ffffffe7399cf339ced6b4e739cf5ab5ad6b5a739cf5ac6b53"),
                (x"fffffce739b5a739ced6b5adad5a739ced39ce739cf5ad4e73"),
                (x"fff39ce6739da79ce6d6b4e69d5ad69a6739cf53d6b58d6b53"),
                (x"fff39ce6739da73b5ad39eb499da73d6a739ce7ac63589eb5a"),
                (x"fff39ce739cdad9b5ad34a53ad5b5ac4e694e31ac635ad6b5a"),
                (x"fff39ce739cdad9b5ad34a53ad5b5ac4e694e31ac635ad6b5a"),
                (x"fff39ce739ce733b5ad6c25294ce73d6b494a53ad6b5a4e318"),
                (x"ffd8cce739ce733b5ad34e3094eb5a9ce78c2529c63094a53a"),
                (x"fff39ce739ce673b5ada4a5294a5294ea739e1294a75ac6b5a"),
                (x"ffd8cce739ce739ce733d6b58c2529d6b139da78d6a769ce73"),
                (x"ffd8cce739ce739ce733d6b58c2529d6b139da78d6a769ce73"),
                (x"fffdece739ce739ce6d6b5ad39cf5a9ea76b5ad3b5a73b5ad3"),
                (x"fffffce739ce6799ce73d4e76b5ad6b5ad6b5ad6b5a7a9ce73"),
                (x"ffffffe673b67369ce799dad3cdad6b5ad6b4e739ced3b4e73"),
                (x"ffffffe739cce79ce739cce79ce739b5ad6b6733b5ad6b4e6c"),
                (x"ffffffe739cce79ce739cce79ce739b5ad6b6733b5ad6b4e6c"),
                (x"ffffffe739ce679ce7399e739cced6b5ad9ce7399ce73cce79"),
                (x"ffffffff39ce739ce739ce739cdad6b5b39cb3d9ce739ce739"),
                (x"fffffffffff3339ce739ce739ce6739e739cfbd9ce72cce739"),
                (x"fffffffffffffec63339ce739ce739ce73ef3bde6318cf318c"),
                (x"fffffffffffffec63339ce739ce739ce73ef3bde6318cf318c"),
                (x"fffffffffffffff6332cce739fff39ce59ffffdef79cef39ce"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffff7fff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_1_0
                (x"ffffffffffffffffffffffffffeb5a9ea739cf3fffffffffff"),
                (x"fffffffffffffffffff99ce79633decfffffffffffffffffff"),
                (x"ffffffffffffffffff39b5ad3ce739ce7fffffffffffffffff"),
                (x"ffffffffffffffffff39b5ad3ce739ce7fffffffffffffffff"),
                (x"ffffffffffffbd9ce673b5ad6b6739ce72c63bffffffffffff"),
                (x"fffffffffffb3d9ce6d6b5ad6b4e73ce739cb3bfffffffffff"),
                (x"ffffffffffeb339ce6739dad39dad6b6739ce59effffffffff"),
                (x"ffffffffffeb339ce6739dad39dad6b6739ce59effffffffff"),
                (x"ffffffff39cb339ce673b5ad69dad6b5b39ce7399cffffffff"),
                (x"ffffffb273b67399ceda9dad6b5ad6b5b339dad69cd9ffffff"),
                (x"ffffffe739b4ed69ce7ad5ad69ce739ce739dad69cf3dfffff"),
                (x"ffffffe7399dad6d6b58d4e739a75ac27139dad3ce72cf7fff"),
                (x"fffffce6739dad34a53ad6b53d25294eb5ad4ed69cf3967fff"),
                (x"fffffce6739dad34a53ad6b53d25294eb5ad4ed69cf3967fff"),
                (x"ffd8ccda73cceda4a5389ce7a4a529d5a78c6ad69cf39fffff"),
                (x"fff39cda73ce6d3d6b49d63094a75ad5a78c6ad69ced6fffff"),
                (x"fff39ce6739cf5ad6b094a5284a718c69294ead6b5ad3cffff"),
                (x"fff39ce673b4d29d69384a5284e1294a758c4ed6b5ad9cffff"),
                (x"fff39ce673b4d29d69384a5284e1294a758c4ed6b5ad9cffff"),
                (x"fff39cced69cf094a529c2528425294e276b5ad6b5a79cffff"),
                (x"fff39cdad6b4f094a5384a52842129c2756b4ed69cf39cffff"),
                (x"fff39ce6d6b5b494a5294210842129c253ad6356b5b39cffff"),
                (x"fff39cce73d6a7a9cf494210842129c271ad6933b5b2c67fff"),
                (x"fff39cce73d6a7a9cf494210842129c271ad6933b5b2c67fff"),
                (x"fff39cdb5a9dad6b5b494e30842129c2676b4f5ab5b3dfffff"),
                (x"fff39ccf5ad4e7ac61294a52842129c27539ced3b5a79fffff"),
                (x"fff39ccf18c4f494a5384a108425294a538c6ad6b5a7967fff"),
                (x"fff39cce739cd294a5384a528425084613ad4ed69cf39cffff"),
                (x"fff39cce739cd294a5384a528425084613ad4ed69cf39cffff"),
                (x"fffffce673b4d294a5294a528421084271ad4f39ce739fffff"),
                (x"fffff667399da7a4a52942108421084e3139ce7963199fffff"),
                (x"ffd8cce673b5ad6d69384a108421294a7139ead3ce599cffff"),
                (x"fff39ce673b5ad3d692942108421294a756b4f53ce72c67fff"),
                (x"fff39ce673b5ad3d692942108421294a756b4f53ce72c67fff"),
                (x"fff39cced6b5ad3c612942108421294a676b4d3ace59e67fff"),
                (x"fff39ce6d6b5ad6d692842108421294a676b5a739cd9eeffff"),
                (x"fff39ce673b5ad69cd294a108421084a756b5b499cf2ef7fff"),
                (x"fff39ce739b5ad6b5b4942108421084a756b5a7a9cf2c67fff"),
                (x"fff39ce739b5ad6b5b4942108421084a756b5a7a9cf2c67fff"),
                (x"fffffcb18ccdad69cf494a5294210842676b5a76ce59ffffff"),

                -- 7_explosion_1_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fe739ce73967ff9ce739ce739ce739cb3fffffffffffffffff"),
                (x"fe739ce73967ff9ce739ce739ce739cb3fffffffffffffffff"),
                (x"ce739ce739cb339ce739ce739ce739ce73ffffffffffffffff"),
                (x"66739ccf39ce7339ce769e7369e739b5b39ce59fffffffffff"),
                (x"66673b5a739e673c635a9dad6b4e739ce79ce679ffffffffff"),
                (x"66673b5a739e673c635a9dad6b4e739ce79ce679ffffffffff"),
                (x"cdad6b5ad6b4ed3c6353d5ad69da73ce6739dad9ef7fffffff"),
                (x"b5ad6b5ad6b5a739ce76d5ad39ce73cced6b4f2c6319efffff"),
                (x"b5ad6b5ad6b4d29d6a769eb58c275ab5ad6b5b39ce7defffff"),
                (x"b5ad6b4e73b69294a756d25294a75a9ea76b5b39ce739fffff"),
                (x"9da73d635ad25294a7169a5294eb5ad253ad4e79ce739fffff"),
                (x"9da73d635ad25294a7169a5294eb5ad253ad4e79ce739fffff"),
                (x"d69294a5294a5294a53ad25294a718d253ad4ed39ced3cffff"),
                (x"4a52942529c2538c61294a5384e1294e358c6b539ced3ce73f"),
                (x"4a129421084a1294a52942109c2529d4f5ad6a769ced6b4e7f"),
                (x"4a108421084212942138421094a529c4f539dad6b5ad6b4e7f"),
                (x"4a108421084212942138421094a529c4f539dad6b5ad6b4e7f"),
                (x"4a10842108421084210842108421084ea739dad69ced69e73f"),
                (x"4210842108421084210842108425294a7539ced39ced6cb19f"),
                (x"4210842108421094a508421084e1294a5294ced6b5a79cb19a"),
                (x"421084a5294a1084a5294a5294a718d253ad4ed6b5a79cfbda"),
                (x"421084a5294a1084a5294a5294a718d253ad4ed6b5a79cfbda"),
                (x"425294a5294a5084a718c63184a718d6938c4ed6b5b39ce733"),
                (x"4a5294a5294e1384a5294a529c275ab5b494ced6ce739cfffa"),
                (x"9eb5a9cf5ac63094a753c253a9e9299cf58c4f39ce739ffff3"),
                (x"b5ad6b5ad69cf5ac6276d6b56b6129c63539ce79ce72cffff3"),
                (x"b5ad6b5ad69cf5ac6276d6b56b6129c63539ce79ce72cffff3"),
                (x"b5ad6b4e73d4e73d6a73d6313b4f5ad6a76b5ad9ce58effff3"),
                (x"9cf5a9a75ab4f36b5ada4eb56b5ad6b5ad6b5ad9633bfffff9"),
                (x"b69299ea739e736b5a7a9dad6b5ad6b5ad39dad9f7bfffffff"),
                (x"cce739e739cb333b5ad6b5ad3b5ad69ce79cce73ffffffffff"),
                (x"cce739e739cb333b5ad6b5ad3b5ad69ce79cce73ffffffffff"),
                (x"6673963339633399ce79ce7399dad6b6739ce59fffffffffff"),
                (x"fb1cef798cce739ce73d66739ce673b672c677ffffffffffff"),
                (x"fb3deeb18ccfff9633ff66739ce739ffd9ef7fffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_1_2
                (x"ffffffb339b4ed69cd28421084a5294ea76b5ad963199fffff"),
                (x"ffd8c66673d4ed6d692942108421084ead6b5ad6ce739cffff"),
                (x"fffde766734ead6d692942108421294a676b5ad69cf39cffff"),
                (x"fffde766734ead6d692942108421294a676b5ad69cf39cffff"),
                (x"fffbdf32739ced69cd294a1084210842756b5ad6b5b39cffff"),
                (x"ffd8cf3339d26769cd294a108421084a7139dad6b5a79cffff"),
                (x"ffd8c667399ea76d69294a108421084a7539dad69cf39cffff"),
                (x"ffd8c667399ea76d69294a108421084a7539dad69cf39cffff"),
                (x"fff39cb3399db53c61294a10842129c2756b5ad69cf3967fff"),
                (x"fffffcb18ccce73c630942108421084a53ad4ed3ce72cfffff"),
                (x"fffffce739ce67ac612842108425294a5294a6769cf39fffff"),
                (x"fff39ce673b5a7a4a7084252842529c25294a6739ce79cffff"),
                (x"ffd8ccced6b5b584a5294a52842129c25294ea78c6279cffff"),
                (x"ffd8ccced6b5b584a5294a52842129c25294ea78c6279cffff"),
                (x"fffffcced69da73d69384a108425294a71ad4e7ad6a79cffff"),
                (x"fffffee6d6d6a769cd384a108461294ead6b5ad3d6ad9cffff"),
                (x"ffd8c666d69a75ac61384a108421084ea7ad4f5a9ce79cffff"),
                (x"fff39ce6d6b6b1a4a5384a108421084a5294ead6b5b39cffff"),
                (x"fff39ce6d6b6b1a4a5384a108421084a5294ead6b5b39cffff"),
                (x"fff39ce673b5a76d69384a10842529c25294e276b5ad9cffff"),
                (x"fff39cced6b5ad69cf094a528427184a5294e273b5a79cffff"),
                (x"fff39cdad6b5a78d69294e30942529c27494a6769cf39cffff"),
                (x"fff399dad6b5b494a758c2529425294e35ad6a739cf39cffff"),
                (x"fff399dad6b5b494a758c2529425294e35ad6a739cf39cffff"),
                (x"fffffb5a73b5b589cedad25294e35a4eb539db399ced9cffff"),
                (x"fffffce673b5b589ceda4a529d4e73c253ad5a799ced967fff"),
                (x"ffd8cce673b5a7ad6b494a53a9eb5ad25339dad39cf39fffff"),
                (x"fffde667399dad3c6138d25339cf5ac6b56b5ad3ce73ffffff"),
                (x"fffde667399dad3c6138d25339cf5ac6b56b5ad3ce73ffffff"),
                (x"fffffee673b5ad39ce739ce73b5b5ad4e76b5a76ce73ffffff"),
                (x"ffffffb273b5ad3ce6d6b5ad6b5a73d5a79ce7369cd9ffffff"),
                (x"fffffffe73ce739ce6d6b5ad3b5ad69cf39ce599ce7fffffff"),
                (x"fffffffffff3339ce736b5ad39da739cf39ce59dffffffffff"),
                (x"fffffffffff3339ce736b5ad39da739cf39ce59dffffffffff"),
                (x"ffffffffffff599ce7399ce76b5ad6b5b39cf99fffffffffff"),
                (x"ffffffffffffdccce739ce736b5ad69cf39cfbdfffffffffff"),
                (x"ffffffffffffffffff39ce7399dad6ce7fffffffffffffffff"),
                (x"fffffffffffffffffff9f318ccce73cfffffffffffffffffff"),
                (x"fffffffffffffffffff9f318ccce73cfffffffffffffffffff"),
                (x"fffffffffffe6739cf53d6b5ffffffffffffffffffffffffff"),

                -- 7_explosion_1_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffe633ffce739ce58cffd99cfff96319df319f"),
                (x"ffffffffffffffe633ffce739ce58cffd99cfff96319df319f"),
                (x"fffffffffffffacce7369e739ce58cee739ce739633de7319f"),
                (x"fffffffffffb339ce736b5ad3ce739cce79ce58cce58cce72c"),
                (x"ffffffffff9ce799ce73b5ad69dad6b5ad39e599ce7339ce79"),
                (x"ffffffffff9ce799ce73b5ad69dad6b5ad39e599ce7339ce79"),
                (x"ffffffffdecdad3b5ad6b5ad6b5a73d4ed6b67339cf534eb56"),
                (x"cffffff58ccdad6b5ad6b5ad6b6929d5ad6b6676d6933d4e73"),
                (x"9ffff73339cdad69cf5ad4e769e35a9cf539ce7a9ce76b5ad6"),
                (x"9ffff66739cce73d6b184e316b6b5ab4f1ad6a73b5ad6b5ad6"),
                (x"9ffffce739ce678d6a734eb53d27189e9294e318d6a73d6b53"),
                (x"9ffffce739ce678d6a734eb53d27189e9294e318d6a73d6b53"),
                (x"d7f39ce739b5a69d6ad6d25384a5294a538c27094a5294a529"),
                (x"9e739ce6d6b5a784a75ac2529c6318c6128421294a5294a528"),
                (x"d7b39cced6b5a7a4a53ac25294a5294a528421094a52942108"),
                (x"d3339cced6b5a694a5294e30942108421294a1084210842108"),
                (x"d3339cced6b5a694a5294e30942108421294a1084210842108"),
                (x"fb339b5a739da73d69294a5284210842108421084210842108"),
                (x"fe673b5a73b5ad39cf49421084210842108421084210842109"),
                (x"fced6b5ad6b5ad3d6a784a5294a108c25094a5084210842109"),
                (x"fced6b5a73b4f5ad6a7a4a5384a1084a5294a509421084a109"),
                (x"fced6b5a73b4f5ad6a7a4a5384a1084a5294a509421084a109"),
                (x"fe7399da739eb58d6b094e309c25294a718c25384a5284a529"),
                (x"fff399da739da7a4a53ac25294a75ad25294a5294a5294eb5a"),
                (x"fffffce739cce7a4a53ad6b494a673b61294a53ad6b1a9dad3"),
                (x"fffffce739ce6d69cf53d25294a75ab69294a7569ce76b5ad6"),
                (x"fffffce739ce6d69cf53d25294a75ab69294a7569ce76b5ad6"),
                (x"ffffff7b39ce6d6b5ad6d2538c6a73b4f494a676b5ad6b5ad6"),
                (x"ffffff318c66676b5a799ce739db5ab4e739ced6b5ad6b5ad6"),
                (x"ffffffffbdcdad39cf399dad3b5b5a9eb139da76b5ad6b5ad9"),
                (x"ffffffffffccf399ce739ce76b5a73d6b139cf339ced69e72c"),
                (x"ffffffffffccf399ce739ce76b5a73d6b139cf339ced69e72c"),
                (x"fffffffffffb339ce6d6ce733b6673b4e739e739ce679ce72c"),
                (x"fffffffffffffffce739ce739ce739ce739ce599ce739ce739"),
                (x"fffffffffffffffffd99ce739ce739ce739cffecce739ce73f"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_2_0
                (x"ffffffffffffffffffffce73e6331867bfffffffffffffffff"),
                (x"ffffffffffffffffffecce7399dad6cb19ffffffffffffffff"),
                (x"fffffffffffffee6318cce7399dad69e739cfbdfffffffffff"),
                (x"fffffffffffffee6318cce7399dad69e739cfbdfffffffffff"),
                (x"fffffffffffffccce679ce7399dad6b5a79cb199ffffffffff"),
                (x"ffffffffffffbd99ced6b5ad6b5a739da79ce739f7bfffffff"),
                (x"ffffffffff77b39b5ad69ce73b5a73c4ed6b67396319ffffff"),
                (x"ffffffffff77b39b5ad69ce73b5a73c4ed6b67396319ffffff"),
                (x"fffff9e58c76739b5ad69dad39cf18423139dad6b598cfffff"),
                (x"ffffff333966679b5ada9dadac612942316b5ad6b5a6cf7fff"),
                (x"fffffff58cf32d39cf49c6b584a5294213ad5ad69cf3d77bdf"),
                (x"ffffffe739666d6b5a694a529c252942118c4ed69cf2c67bdf"),
                (x"fffff666d69ced6b5929421084a5084211ad4ed6b5b3967bdf"),
                (x"fffff666d69ced6b5929421084a5084211ad4ed6b5b3967bdf"),
                (x"fffffce6d6b5ad69cd084210842108421094a756b5a79cb19f"),
                (x"fffffcce73b5ad69cd284a1084210842118c2756b5ad39e73f"),
                (x"fffffccf399ce769cd284252842108425294a7539cf33ce73f"),
                (x"fffffce739cce73d69284a109421084a5084275ad6b59ce73f"),
                (x"fffffce739cce73d69284a109421084a5084275ad6b59ce73f"),
                (x"fff39ce739cdada4a7184a10845d08425084267ad6a73ce73f"),
                (x"fb339ce7399cf584a52942108b86f74210844ed39ced967bdf"),
                (x"fe7399e6739e929421184210845c21ba1294ea739ce6c77bdf"),
                (x"fe739b5ad6b6929421294211bbdc21ba1094ea739ced977bdf"),
                (x"fe739b5ad6b6929421294211bbdc21ba1094ea739ced977bdf"),
                (x"ff7bdcce739ce7a4a50842101ba37bda1294e1299ce7967bdf"),
                (x"fffde64d294ea7a4210842101ba108427094a1099ced9639df"),
                (x"fffff6675ad6b5a4a50842117da10842108421099ce79efbdf"),
                (x"fffff666d6b5ad8421084210842108421084213a9cf3d77fff"),
                (x"fffff666d6b5ad8421084210842108421084213a9cf3d77fff"),
                (x"fffde666d69ea69421084210846f7b421294a3099cd8ef7fff"),
                (x"ffbbdcdad69e9284210842108d8421ba13ad635a9cf39f7bdf"),
                (x"ff98ccced6b4f094210845efbb84210a138c275a9ced9f7bdf"),
                (x"ffbde666d6b4d294a50846f770def70dd139ce699ced3cfbdf"),
                (x"ffbde666d6b4d294a50846f770def70dd139ce699ced3cfbdf"),
                (x"fe739cdad6b4d294a50845ef7ba2f70ed18c6a73b5b39cb19f"),
                (x"fff39ce673d4f494a50846f7708421ba138c2716b5a79ce73f"),
                (x"fffbd67b399db49c610846f77bdef70dd139ce76b5a79ce73f"),
                (x"fbbdece673d4f494a70945ef708421bed094eb56b5a79cb19f"),
                (x"fbbdece673d4f494a70945ef708421bed094eb56b5a79cb19f"),
                (x"fb33967b399db49c630946f7bb86f7da10842676b5a79cb9df"),

                -- 7_explosion_2_1
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"63bfffe7def7bffffffdce72cfffffffffffffffffffffffff"),
                (x"cfbbdce7de677dffffddce739cffffffffffffffffffffffff"),
                (x"cfbbdce7de677dffffddce739cffffffffffffffffffffffff"),
                (x"6658cce58cce58c63199b4e79ce739ce59ffffd3ffffffffff"),
                (x"f67decdb399db39ce673b6739ce6739e739cf599ffffffffff"),
                (x"ccf399dad6b5ad6d6933b4e79ce7399dad9cb32cffffffffff"),
                (x"ccf399dad6b5ad6d6933b4e79ce7399dad9cb32cffffffffff"),
                (x"9ea73d5ad6b4e76d6933b4e73ce673b5a6c6798e73bfffffff"),
                (x"b4ed69ce739eb56d6b53d6b53b4e73b5a79cb339f7bdffffff"),
                (x"d6b5ad2529c2676d6a734a53ab4e73b5ad6b5a79ce7defffff"),
                (x"4a5294a5294a138d6b5a4a538d4ed6b5ad6b4f39ce72c77fff"),
                (x"c27184a529421084a509421094ea739ced6b4ed6b5a7967fff"),
                (x"c27184a529421084a509421094ea739ced6b4ed6b5a7967fff"),
                (x"c61084210842108421084a109c25294a1339ead6b5ad367fff"),
                (x"4a5084210842108421084e309c2108421294a756b5ad96319f"),
                (x"42108421084210842108421084a5084a1094e2739ced9ce739"),
                (x"ddf7bddf7bba108421084210842129421094ead69ced9ce739"),
                (x"ddf7bddf7bba108421084210842129421094ead69ced9ce739"),
                (x"ddef7bdef7da108bdc21da10842508421094e3539ced9ce73e"),
                (x"b86f70dc21bed08deef7ba1174210842138c2713b5ad39ce6c"),
                (x"086f70a2f70876842108bdee1ba108421294a713b5ad6b5acc"),
                (x"b86f70def7087684211b0843742108421094a5389ce76b5ad8"),
                (x"b86f70def7087684211b0843742108421094a5389ce76b5ad8"),
                (x"ddc21b84210dd084211bbdee8425084210842108c62769e72c"),
                (x"46ef746ef74210842128421084a52942108421089ced6cb19e"),
                (x"421084a1084a5284230942528421294210842718b5a73cb19f"),
                (x"42673c6273c6928421294a52842129c2758c6ad3b5b39cffff"),
                (x"42673c6273c6928421294a52842129c2758c6ad3b5b39cffff"),
                (x"4ea734ea734e10842118d6b534a5294a6739dad6ce72cf7fff"),
                (x"9ea73c4e73d6b09421099ce769eb5ad6ad6b5ad6ce72cf7fff"),
                (x"b5ad6b4d29d693a4a5299ce73d6a73b5ad6b5ad6ce739fffff"),
                (x"b5ad6b5a739ce739ce739ce73d6a73b5ad39ced6633dffffff"),
                (x"b5ad6b5a739ce739ce739ce73d6a73b5ad39ced6633dffffff"),
                (x"9ce739e6d6b65999ced3b4e769eb39b4f39ce66c633fffffff"),
                (x"ce739ce673ce5ddce739cb1999e6739e72c6758cffffffffff"),
                (x"ce739ce739f7bceef58c739ccce7399e58c63bdfffffffffff"),
                (x"73339cb3def7bfff79def7bdece739cb3def7bffffffffffff"),
                (x"73339cb3def7bfff79def7bdece739cb3def7bffffffffffff"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_2_2
                (x"fbb39cced6b4d284211bb8437ded084e3094ead3ce7cccb19f"),
                (x"fb339cced6b6b494237708421bdd084e1294ea7a9cf39f39df"),
                (x"fe739cced6b4e73422e1bdef7bed08423094ead3ce7cceffff"),
                (x"fe739cced6b4e73422e1bdef7bed08423094ead3ce7cceffff"),
                (x"fe739cced6b61384a51708421bed08421294ea7a9cf39cffff"),
                (x"fb339ce6d69cf5842361ba117bdd08421294a676b5ad9ce73f"),
                (x"ffb399da734ce73422e1bdee1bed08421294a676b5b2cf7bdf"),
                (x"ffb399da734ce73422e1bdee1bed08421294a676b5b2cf7bdf"),
                (x"ffbdecda73d69384a50108437ddd08421094e276b5a7967bdf"),
                (x"ffbdece673d6b1a4a5170843b421084210842753b5ad9efbdf"),
                (x"fffde732734e1094a508def6842108421094cf53b5b2cf7fff"),
                (x"ffdceee673d250842108421084210842118c5ad6b5b2cfffff"),
                (x"ffbbdcce734a108421084211bba1084213ad6b5ad6b2cfffff"),
                (x"ffbbdcce734a108421084211bba1084213ad6b5ad6b2cfffff"),
                (x"fb98ccda734a109c6128421170a1084211ad4f494a66cf7fff"),
                (x"ff98ccce734a7094a51bda1170a1084213ad4e739ce79ef7bf"),
                (x"ff9cecda739cf49421170def7da1084a5094a756b5ad6ce73f"),
                (x"ff9ce64e739cf494a5170dee842108c21094a7539cf33ce73f"),
                (x"ff9ce64e739cf494a5170dee842108c21094a7539cf33ce73f"),
                (x"ff98ccda739da6842108b8437421084a538c6a73ce739cb19f"),
                (x"fe7399cf5ad4d284212845ee842129c613ad5ad9ce739cffff"),
                (x"fe739ceb5ad692842129421084a129427539ce79ce739fffff"),
                (x"fe7399e6739e9294a528421084250842676b4e73ce679fffff"),
                (x"fe7399e6739e9294a528421084250842676b4e73ce679fffff"),
                (x"fe6739dad6b693842108421084212942676b5ad69ce79fffff"),
                (x"fb339cced6b692942108421084210842276b5ad6b5b39fffff"),
                (x"ff98cce6d6b5a7a4210842529421084a6d6b5a73b5b2cfffff"),
                (x"ff98c66673b5a78421084a5384a5294ced6b5b2cce73ffffff"),
                (x"ff98c66673b5a78421084a5384a5294ced6b5b2cce73ffffff"),
                (x"ff9ceee673b5ada4a5084a529c6b184ea739d99e633bffffff"),
                (x"fffde64ed6b5ad6c61084e318d5a73d5ad9ccf2cce59efffff"),
                (x"fffff632d6b5ad3c6108c4e739da73b5ad9ce72e63333fffff"),
                (x"ffffffb18cce736b5a789dad69ce73b5ad9ce7ceffffffffff"),
                (x"ffffffb18cce736b5a789dad69ce73b5ad9ce7ceffffffffff"),
                (x"ffffffffdece7399ced39dad6b5ad6b5a79cfbdfffffffffff"),
                (x"ffffffffffcb1999ced6b5ad3ce739ccf2c67bffffffffffff"),
                (x"ffffffffffffbd9ce733b5ad3ce7396318e77fffffffffffff"),
                (x"fffffffffffffff63199b5ad3ce73967ffffffffffffffffff"),
                (x"fffffffffffffff63199b5ad3ce73967ffffffffffffffffff"),
                (x"ffffffffffffffffffccc318cf6739ffffffffffffffffffff"),

                -- 7_explosion_2_3
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffdef7999ce739f7bdef3bdffffdef7999cb18e"),
                (x"ffffffffffff9cc63333ce739639ce633ae77bdece739ce739"),
                (x"ffffffffffff9cc63333ce739639ce633ae77bdece739ce739"),
                (x"ffffffffff633acce7339e733cb339ce73debb399cf39ce739"),
                (x"fffffffd8c64f39ce676ceb53b4ed69da79cb336b5b339ce73"),
                (x"fffffff98cb5a73b5ad69eb5a9ce739ce739ce739ced6b5ad6"),
                (x"fffffff98cb5a73b5ad69eb5a9ce739ce739ce739ced6b5ad6"),
                (x"fffffce739b5ad6b5ad69eb5a9ce734a53ad275a4a676b5ad6"),
                (x"fffde66739b5ad6b5b5ad6b53b4e734a1094e35a9ce789eb53"),
                (x"fffde66739b5ad39cd294a5299eb5ac2108423099cf499eb49"),
                (x"fff39ce6d69db58d69384a108425294a508427589cf189a528"),
                (x"fb3399ced6c6128421084a108425084e108425294210942108"),
                (x"fb3399ced6c6128421084a108425084e108425294210942108"),
                (x"f3339b5a7342108421084a529421084250842108bdf68bef68"),
                (x"66673b4f1842108421084252845ef7da108422e1084370defb"),
                (x"c5ad6b4e73c25294210842108b8421da10846c21bdee1b8437"),
                (x"65ad6b5ad69e1294a508421170def74210846c21bdd01b8421"),
                (x"65ad6b5ad69e1294a508421170def74210846c21bdd01b8421"),
                (x"64e739dad69e1384a50842108ba2f7bdf6842377086e1b8437"),
                (x"f6739cda739eb0942108425284237b086e84211bbdef7bdefb"),
                (x"ce739cda73b5b49421084a108421084210842117deefbddefb"),
                (x"ce739cda739cf0942109425294210842108421084210842108"),
                (x"ce739cda739cf0942109425294210842108421084210842108"),
                (x"fb18ccdad6b69294a508421184e12942108421084210842529"),
                (x"ffd8c9dad6b5b534a5094a5384a12942108421084210846318"),
                (x"ffd8ccced6b5a76b5a739eb494a1084a128421084a529c2538"),
                (x"ffdce66739ce676b5ad6b4e7ac2529d6b58c25094a5294a529"),
                (x"ffdce66739ce676b5ad6b4e7ac2529d6b58c25094a5294a529"),
                (x"ffffff7b39cced6b5ad69ce76d25299cf56b4d384a53ad6b5a"),
                (x"fffffffbdece5999ced69ce769eb5a9eb56b6b539ce73b4e76"),
                (x"fffffffdce733cc9ced69e7399ced69a756b4e76b5ada9eb53"),
                (x"ffffffffff66599b5ad3ce739cced69a756b5ad6b5ad3cce79"),
                (x"ffffffffff66599b5ad3ce739cced69a756b5ad6b5ad3cce79"),
                (x"ffffffffffcb3b9ce7339e739ce6d69cf39ce6d3ce6d9f673e"),
                (x"ffffffffff9fbff63339ce739cced6cb18c63339633396672c"),
                (x"ffffffffffffffffffffffff9ce739efbffffbacf7b39efbd9"),
                (x"fffffffffffffffffffffffff66739efffffffdef7b3ffb9cc"),
                (x"fffffffffffffffffffffffff66739efffffffdef7b3ffb9cc"),
                (x"ffffffffffffffffffffffffffffffffffffffffffffffffff"),

                -- 7_explosion_3_0
                (x"cfffffffffffffdce739cce739e6734a53ad7fffffffffffff"),
                (x"ffffffffffffff9ce6739dad6b66739cf4c67fffffffffffff"),
                (x"ffffffffffb5b39b5ad6b5ad6b5a73ce72c633ffffffffffff"),
                (x"ffffffffffb5b39b5ad6b5ad6b5a73ce72c633ffffffffffff"),
                (x"fffffffed6b5ad39ced6b5ad6b5a739ced39ce7fffffffffff"),
                (x"ffffffdad6b4f49d6ad69ce769dad69db5ad599effffffffff"),
                (x"ffffffcf5a9cd29d6a769ce76d6b5a9da78c4ecc633fffffff"),
                (x"ffffffcf5a9cd29d6a769ce76d6b5a9da78c4ecc633fffffff"),
                (x"ffffffe929d69384a7099dad3c2718b5b494ead9ce5dffffff"),
                (x"fffffb6929c210842129c4e784a5299db494e273633d6fffff"),
                (x"fff39b6929c250842109c6b494a108425294e13ace6d667fff"),
                (x"ffe739e1294a5094a5084a52942108421094a533b5ad6cffff"),
                (x"ffd8cce9294a1094a5284210942108421294a2769cf2c67fff"),
                (x"ffd8cce9294a1094a5284210942108421294a2769cf2c67fff"),
                (x"fffdeccf5a4a5084a52842108421084210842756b5b3967fff"),
                (x"fffbdcdb5a4a1094a508421084237b4210842756b5ad6cffff"),
                (x"ffbde9db5a4a508421084210846f7b4210842356b5ad6cf7bf"),
                (x"f33bdb5a73c252842117bef6845f7b4210842118d6b539b18c"),
                (x"f33bdb5a73c252842117bef6845f7b4210842118d6b539b18c"),
                (x"f673965ad6b6929421170dee10def742108421084a53ad6739"),
                (x"ce7399ced6b6908421170def7b86f742108421084a53a9e739"),
                (x"cb3def6739b690842361b8437dec21da108421084a7139e739"),
                (x"fb1cef3339b4d08dec21bdef70a2f7ba1094a109d6a6c6673f"),
                (x"fb1cef3339b4d08dec21bdef70a2f7ba1094a109d6a6c6673f"),
                (x"fffdef32734a508deef74211708421da1294a5299cede77fff"),
                (x"fffde665294213842368ddef708421da108421099ceccf7fff"),
                (x"ffdceecf184212942117bdee10dc21da10842108c6273f7bdf"),
                (x"ffd8cccd0842108def7708421bdc210dd08421084a756cb18c"),
                (x"ffd8cccd0842108def7708421bdc210dd08421084a756cb18c"),
                (x"ffed6b4d29421084236108437ded0845efbda108423569e739"),
                (x"ffed6b5b5a4210842117bdef70dd08b84210ed08423569e739"),
                (x"732d69cf5a4a1084a51bbdee1086f7b8768421084227367bde"),
                (x"67a73d6129425284a517084210df7bba108421084a6d9f7bdf"),
                (x"67a73d6129425284a517084210df7bba108421084a6d9f7bdf"),
                (x"cb3399a71842528c6137b8421086f7da1084210842279f7fff"),
                (x"ce7399ea734a1384a51b45ee1084210ed08421294a66c77fff"),
                (x"ce6739da734a1094210845ee108421ba1084211a9ce6cf7fff"),
                (x"fe673b4f184a1084210846f77084210dd084211ab5acc77fff"),
                (x"fe673b4f184a1084210846f77084210dd084211ab5acc77fff"),
                (x"fff5a9e929d21084210842117b8421ba10842113b5acc77fff"),

                -- 7_explosion_3_1
                (x"fff39ce58c77fffffffffe739f7bfffffffffffffffffffff9"),
                (x"fe739cb3de67ffffffff63199cb3deffffffffffffffffffff"),
                (x"d4e73ce673b5acc73bde77bd9cf7deef9939e7ffffffffffff"),
                (x"d4e73ce673b5acc73bde77bd9cf7deef9939e7ffffffffffff"),
                (x"9da739cf5a9dad9ef59ef7bd365a73ce7339dadfffffffffff"),
                (x"d4ed6d27189da739cf2c66733b5ad6b4f58c6b5a9cedffffff"),
                (x"4e2739e129d6928c6133ce736b4f5ad69294a529d6ad6fffff"),
                (x"4e2739e129d6928c6133ce736b4f5ad69294a529d6ad6fffff"),
                (x"d25294a1084a10842109b5ad6b61294a5294e31a9ced6b7fff"),
                (x"421084252942108421099eb5ad2529425094a51a9ce76b7fff"),
                (x"421084a529421084a528421084a50842108421094a756cffff"),
                (x"42129c2108421084a708421084a1084a1294a1184a533ce73d"),
                (x"421084e1294a11b4211bda108421084a5294a109d6b53b6739"),
                (x"421084e1294a11b4211bda108421084a5294a109d6b53b6739"),
                (x"42108425084237b423770ef684210842528421389ced6b4e79"),
                (x"42108ddef7ddc37bdd1708437bdd084210842529b5ad6b4e79"),
                (x"4210845c21bdc21bdf68bdee10dd08421094e3139ce76b4e79"),
                (x"46ef7b8421bdc21bdee8b8437bed08421094ea769ce76b5ad3"),
                (x"46ef7b8421bdc21bdee8b8437bed08421094ea769ce76b5ad3"),
                (x"bdc21084210dee1086f7bdef70a108421294a713b5ad6b5ad3"),
                (x"b84210842108777084210ef770a1084210842538d6a76b5ad3"),
                (x"08421086f70df77bdc2146f61bdf7b4210842129d6ad6b6739"),
                (x"084210df7bba10108421b8437bef7bda10842138d6ad39ce73"),
                (x"084210df7bba10108421b8437bef7bda10842138d6ad39ce73"),
                (x"b86f70eef7bdd01def7bbef684210842108422769ce73cce69"),
                (x"45d08da108086f742108421084210842108426d6b5ad3cce69"),
                (x"4210842108d86e8421094210842108421284275a9cf56ceb49"),
                (x"421084210840768421094a10842108421294a529c63536319a"),
                (x"421084210840768421094a10842108421294a529c63536319a"),
                (x"421084210846d084210942108421084a5094e31a9ced367fff"),
                (x"421084a1084210842109421084235ad6a694a676b5993fffff"),
                (x"9eb5a4a10842108421294a108462d6b5ad39ea79633dffffff"),
                (x"b5a734a12942109c6273d25294ead6b5a76b6599633fffffff"),
                (x"b5a734a12942109c6273d25294ead6b5a76b6599633fffffff"),
                (x"b5a739ced69eb5a9ced69e3094ead6b6736b5bceffffffffff"),
                (x"6318c667399dad69cd9e64e7ad4ed6b6596b5adfffffffffff"),
                (x"73bde77bde64e79f7bce64e73d4f39cb199cb3ffffffffffff"),
                (x"ffffffffdef672cf7bffce739cb3bdffffffffffffffffffff"),
                (x"ffffffffdef672cf7bffce739cb3bdffffffffffffffffffff"),
                (x"fffffffffff672cffffffe739cb3ffffffffffffffffffffff"),

                -- 7_explosion_3_2
                (x"ffdce65ad69a1084211708437ba108421084211a4a753d7fff"),
                (x"ffdce65ad6d2108422e108421bed084210842109c62769e73f"),
                (x"fffde64e73d210842117084210dd08421094a1099ced39e739"),
                (x"fffde64e73d210842117084210dd08421094a1099ced39e739"),
                (x"ffdce64d294a50842361084210dd08da138c25099cf53ce739"),
                (x"fffdeccd08421084211bb8421086f7ba70842528c6133cb199"),
                (x"ffbdecd9294210842117ddee108421ba128425284a71a9fbcc"),
                (x"ffbdecd9294210842117ddee108421ba128425284a71a9fbcc"),
                (x"f798c9cd0842108dec37b84210def7da12842109d6a73b318e"),
                (x"ce673b6908423610843745ee1bdef7ba10842108d6ad6b7fff"),
                (x"ce673b69084211bbdee846f7bb84210ed08421084a676b7fff"),
                (x"63339b692942108422e10def708421bef68421084227967fff"),
                (x"ffbde9cf18421084211b0dee10def7ba1094a508c627d77fff"),
                (x"ffbde9cf18421084211b0dee10def7ba1094a508c627d77fff"),
                (x"fffde65a734a1084211b08421bdf7b46d18c25084a72cf7fff"),
                (x"ffdcef5a734a5294a51b08421ba108bdf68421299cd9ef7fff"),
                (x"fe58c64f5a4a10942117ba101bdef70876842276ce59e7319f"),
                (x"ce6739e129421084211b0ef7bb86f70ed0842356ce73ef3199"),
                (x"ce6739e129421084211b0ef7bb86f70ed0842356ce73ef3199"),
                (x"ce673d25294210842108b8437bdc21ba10842356b5a73ce739"),
                (x"ce75ad25294210842108bdee10dc21ba1094a756b5accce73e"),
                (x"632739eb5ac210842108ddee846ef7ba108425389ced6eb19e"),
                (x"ff739b5ad6b690842108def68421084210842129d6ad3f7bdf"),
                (x"ff739b5ad6b690842108def68421084210842129d6ad3f7bdf"),
                (x"fff39b5ad6b692842108da10842108421294a109d6ad9effff"),
                (x"ffd8cce6d6b69284210842108421084252842129d6a79f7fff"),
                (x"ffd8c66673b4d094a508421084a108425294a1094a75967fff"),
                (x"fff39b5ad69a52942108421084a529421294a1294a7139ffff"),
                (x"fff39b5ad69a52942108421084a529421294a1294a7139ffff"),
                (x"ffd8cb5b39d27094a528421094eb184a108421384a756cffff"),
                (x"fffffb798c9cf09d6ad34a529c4f184a508421184a756fffff"),
                (x"ffffffbb39cdb49d6ad6c25389da734e138c275a4a75ffffff"),
                (x"fffffffd8c65a789ced3d6b5ab4e73b4f494a673d6a7ffffff"),
                (x"fffffffd8c65a789ced3d6b5ab4e73b4f494a673d6a7ffffff"),
                (x"fffffffffff32dad6ad3b5ad3b4e73b5b494ea76b5adffffff"),
                (x"fffffffffffce73b5a739dad6b5ad6b5a739dad6b5bfffffff"),
                (x"ffffffffffffd8cce7399dad6b5ad6b5ad9ce6d6ffffffffff"),
                (x"fffffffffffffecd6a739e736b5a739cf39cffffffffffffff"),
                (x"fffffffffffffecd6a739e736b5a739cf39cffffffffffffff"),
                (x"ffffffffffffffa4a5299e7339cf39ce73defffffffffffff9"),

                -- 7_explosion_3_3
                (x"fffffffffffffffffffffb199ce7fffffec6673effffffffff"),
                (x"ffffffffffffffffffffeb199ce739fffcc6673ef7bfffffff"),
                (x"ffffffffffffd9963199cce7a9cd8c77bd9cce6cf7bcef39ce"),
                (x"ffffffffffffd9963199cce7a9cd8c77bd9cce6cf7bcef39ce"),
                (x"fffffffffffdad663336b4e7ad4d8cf3276b5ad3ce72c6318c"),
                (x"ffffffffff77ad6ce736b6b494e273b5a7ad6b53b5a739dad6"),
                (x"fffffffd8ccb3369ced6b6b494a75a9cf094a1084a5099dad6"),
                (x"fffffffd8ccb3369ced6b6b494a75a9cf094a1084a5099dad6"),
                (x"fffffff98cccf53b5ad6b6308421294a5084210842109d6b53"),
                (x"fffff9b2d6b4d299cf5ad2108421084a108421084210942108"),
                (x"ffd8c9da73d63094212942108421084a108423684210842108"),
                (x"d318c9eb184a5294a50842108421294a10846c284210842108"),
                (x"4eb39b6a73d69284a50842108421084a10845c3b4210842108"),
                (x"4eb39b6a73d69284a50842108421084a10845c3b4210842108"),
                (x"4cf399dad6b592842108421084210842117bdc214211b45ee8"),
                (x"4cf399ce73b4d08421084210846ef7def610a2f7bdf61b8437"),
                (x"9ce739db5ac25084211bdef77b86f7084210a117deee108421"),
                (x"ce6d6b5b5a4a50842108ddef70ed08086f7beee1bdc2108421"),
                (x"ce6d6b5b5a4a50842108ddef70ed08086f7beee1bdc2108421"),
                (x"9dad6b4f5ac25284210842101bec2108437bec210842108437"),
                (x"9dad6b5ad69e1294a50842101bdef7bdc210dee1084210def7"),
                (x"9dad6b4e73b4f494210846f77b86f745ee1086f708437bef68"),
                (x"cced6b4e739e3094210845ee10def746ee1086f7086e842108"),
                (x"cced6b4e739e3094210845ee10def746ee1086f7086e842108"),
                (x"cced6b5ad64a5284210845ef7b8421ba2f7b86fbbdefb42108"),
                (x"cced6b5a73c25084a5284210846c21bed1bded084212842108"),
                (x"ce6d69eb5a4a1094a529421084237bda11bda1094a70942108"),
                (x"ee7399a529c21094a50942109421084612842108421184a108"),
                (x"ee7399a529c21094a50942109421084612842108421184a108"),
                (x"fff39b69294a10842108425294210842528421084a52942108"),
                (x"ffed6b4e73d2129421284a53ad6a734a108421084a52842108"),
                (x"ffed6b5a73d63094a5294e316b5ad64a10842109421094a53a"),
                (x"fffffb5b5a4a5294a75ad4e76b67399a7084275a4a7139e309"),
                (x"fffffb5b5a4a5294a75ad4e76b67399a7084275a4a7139e309"),
                (x"ffffffda73d6b58d6a76b5ad69e58c666739ced3c613ab4e7a"),
                (x"fffffffffffdad3ce7399dacc9fbdef33b9cdad3d6a739dad3"),
                (x"fffffffffffff33633ddf77b9cf9cef79cc65ad69cf399ce7a"),
                (x"fffffffffffffffffffff3199cb18cffffffffecf7999ce73f"),
                (x"fffffffffffffffffffff3199cb18cffffffffecf7999ce73f"),
                (x"cfffffffffffffffffffffbdece7ffffffffffee63339cffff"),

                -- 8_bonus-life
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296736b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6f39ce739ce71ad6b79ce739ce738d6b5ad9cca5"),
                (x"296736b5ad6f39ce739ce71ad6b79ce739ce738d6b5ad9cca5"),
                (x"296736b5b4a4e78c63189ce94a52734a53ad4e74a35ad9cca5"),
                (x"296736b5b4a4e78c63189ce94a52734a53ad4e74a35ad9cca5"),
                (x"29739a52939a528421084a6739cd294211ef6b539d294ce4a5"),
                (x"29739a52939a528421084a6739cd294211ef6b539d294ce4a5"),
                (x"29739a5289484210a1084235ac6108739cb5fbdad5294ce4a5"),
                (x"29739a5289484210a1084235ac6108739cb5fbdad5294ce4a5"),
                (x"29739a5289484210a1084235ac6108739cb5fbdad5294ce4a5"),
                (x"29739a5289484210a108a53bda53bd2108e721094d294ce4a5"),
                (x"29739a5289484210a108a53bda53bd2108e721094d294ce4a5"),
                (x"29739a52894a10845294a508484000ef7a8421094d294ce4a5"),
                (x"29739a52894a10845294a508484000ef7a8421094d294ce4a5"),
                (x"29739a52939a117bd29439ca57bfbda5288421139d294ce4a5"),
                (x"29739a52939a117bd29439ca57bfbda5288421139d294ce4a5"),
                (x"296736b5b4a25284739c319ef73bbde738842534a35ad9cca5"),
                (x"296736b5b4a25284739c319ef73bbde738842534a35ad9cca5"),
                (x"296736b5bce4e78c5294003bdef79ca5298c4e7ce35ad9cca5"),
                (x"296736b5bce4e78c5294003bdef79ca5298c4e7ce35ad9cca5"),
                (x"296736b5bce4e78c5294003bdef79ca5298c4e7ce35ad9cca5"),
                (x"296736b5ad6d2939eb5aa539ce7294d6b539d28d6b5ad9cca5"),
                (x"296736b5ad6d2939eb5aa539ce7294d6b539d28d6b5ad9cca5"),
                (x"296736b5ad6b5b4a5294d69084235aa5294a35ad6b5ad9cca5"),
                (x"296736b5ad6b5b4a5294d69084235aa5294a35ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5adef5294a7bd6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5adef5294a7bd6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b694a51ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b694a51ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b694a51ad6b5ad6b5ad6b5ad9cca5"),
                (x"296739ce739ce739ce739cf39ce6739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739cf39ce6739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 9_bonus-godmod
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739ce739cfbdef6739ce79cce739ce739cca5"),
                (x"296739ce739ce739ce739cfbdef6739ce79cce739ce739cca5"),
                (x"296736b5ad6b5bded294a516b21294a529deb5ad6b5ad9cca5"),
                (x"296736b5ad6b5bded294a516b21294a529deb5ad6b5ad9cca5"),
                (x"296736b5ad6b5bded294a516b21294a529deb5ad6b5ad9cca5"),
                (x"296736b5ad6f38b590841094a5ac425ad64277ad6b5ad9cca5"),
                (x"296736b5ad6f38b590841094a5ac425ad64277ad6b5ad9cca5"),
                (x"296736b5ad6d28a52d6ba50c65acc65294b5d28d6b5ad9cca5"),
                (x"296736b5ad6d28a52d6ba50c65acc65294b5d28d6b5ad9cca5"),
                (x"296736b5ad6f3873a94a3194a5ae9439ceb5884d6b5ad9cca5"),
                (x"296736b5ad6f3873a94a3194a5ae9439ceb5884d6b5ad9cca5"),
                (x"296736b5ad6d28a5294aa514a52a948c62b5f7ad6b5ad9cca5"),
                (x"296736b5ad6d28a5294aa514a52a948c62b5f7ad6b5ad9cca5"),
                (x"296736b5ad6d28a5294aa514a52a948c62b5f7ad6b5ad9cca5"),
                (x"296736b5bded294a739c1084231a94a5294a77ad6b5ad9cca5"),
                (x"296736b5bded294a739c1084231a94a5294a77ad6b5ad9cca5"),
                (x"29673a528b5843def39c5294a8c4e78c634a77ad6b5ad9cca5"),
                (x"29673a528b5843def39c5294a8c4e78c634a77ad6b5ad9cca5"),
                (x"29673a528a52d6b5f7bd39d4a39d6b5ad6a5738d6b5ad9cca5"),
                (x"29673a528a52d6b5f7bd39d4a39d6b5ad6a5738d6b5ad9cca5"),
                (x"29673a529ce294f7ad6b5adcea514a5ad6b5f38d6b5ad9cca5"),
                (x"29673a529ce294f7ad6b5adcea514a5ad6b5f38d6b5ad9cca5"),
                (x"296736b5bce18ca54a520856ba514a5ad718d28d6b5ad9cca5"),
                (x"296736b5bce18ca54a520856ba514a5ad718d28d6b5ad9cca5"),
                (x"296736b5bce18ca54a520856ba514a5ad718d28d6b5ad9cca5"),
                (x"296736b5ad6f3863294a5ad6b1094a529463738d6b5ad9cca5"),
                (x"296736b5ad6f3863294a5ad6b1094a529463738d6b5ad9cca5"),
                (x"296736b5ad6b5bce18c65296ba514a5295ce35ad6b5ad9cca5"),
                (x"296736b5ad6b5bce18c65296ba514a5295ce35ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6d29439d4a31bde318cd6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6d29439d4a31bde318cd6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5bce77bd5294a5ad6b8c63ce35ad6b5ad9cca5"),
                (x"296736b5ad6b5bce77bd5294a5ad6b8c63ce35ad6b5ad9cca5"),
                (x"296736b5ad6b5bce77bd5294a5ad6b8c63ce35ad6b5ad9cca5"),
                (x"296739ce739ce74a739c31842108c6318d4a4e739ce739cca5"),
                (x"296739ce739ce74a739c31842108c6318d4a4e739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 10_bonus-wallhack
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"29673ce739cce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"29673ce739cce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296736b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"294210842422d6b5f39ce73bde739ce739ce77bce739c9cca5"),
                (x"294210842422d6b5f39ce73bde739ce739ce77bce739c9cca5"),
                (x"296736b5ad6fbc21318c18ef718e94631831dee31d294ce4a5"),
                (x"296736b5ad6fbc21318c18ef718e94631831dee31d294ce4a5"),
                (x"297396b5a422d7082d6b5ac6318e946318318c631d294ce4a5"),
                (x"297396b5a422d7082d6b5ac6318e946318318c631d294ce4a5"),
                (x"296736b5ad6fbc63318c6318c632946318c6318c652949cca5"),
                (x"296736b5ad6fbc63318c6318c632946318c6318c652949cca5"),
                (x"296736b5ad6fbc63318c6318c632946318c6318c652949cca5"),
                (x"2967321084214a52c21000000a5294a5294a5294a52949cca5"),
                (x"2967321084214a52c21000000a5294a5294a5294a52949cca5"),
                (x"296736b5ad6fbc6318c61098c18ef718c74a0c652d294ce4a5"),
                (x"296736b5ad6fbc6318c61098c18ef718c74a0c652d294ce4a5"),
                (x"2942121084214ab5ad6b5ad6b18c6318c74a0c631d294ce4a5"),
                (x"2942121084214ab5ad6b5ad6b18c6318c74a0c631d294ce4a5"),
                (x"296736b5ad6fbcc6318c1098c6318c63194a318c652949cca5"),
                (x"296736b5ad6fbcc6318c1098c6318c63194a318c652949cca5"),
                (x"29673210842420000000a5294a5294a5294a5294a52949cca5"),
                (x"29673210842420000000a5294a5294a5294a5294a52949cca5"),
                (x"29673210842420000000a5294a5294a5294a5294a52949cca5"),
                (x"296736b5ad6fbcc60c6318ef718e94631831dee31d2949cca5"),
                (x"296736b5ad6fbcc60c6318ef718e94631831dee31d2949cca5"),
                (x"294212108422d6b5ad6b18c6318e946318318c631d294ce4a5"),
                (x"294212108422d6b5ad6b18c6318e946318318c631d294ce4a5"),
                (x"296736b5ad6ffe6318c6e739ce739ce739ce739ce739c9cca5"),
                (x"296736b5ad6ffe6318c6e739ce739ce739ce739ce739c9cca5"),
                (x"297396b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"297396b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"297396b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad9cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 11_bonus-speed
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296736b5ad6b5ad6b5ada518c6318c6318c6319ce35ad9cca5"),
                (x"296736b5ad6b5ad6b5ada518c6318c6318c6319ce35ad9cca5"),
                (x"296736b5ad6b5ad6b5ada518c6318c6318c6319ce35ad9cca5"),
                (x"296736b5ad6b5ad6b5ade70630856b8420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6b5ade70630856b8420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6f7bd421084a75a8420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6f7bd421084a75a8420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6b5adef6318c6318420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6b5adef6318c6318420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6f39c4a508c62738420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6f39c4a508c62738420a518dce35ad9cca5"),
                (x"296736b5ad6b5ad6f39c4a508c62738420a518dce35ad9cca5"),
                (x"296736b5ad6f394a5294ef6318c6318420a577bce35ad9cca5"),
                (x"296736b5ad6f394a5294ef6318c6318420a577bce35ad9cca5"),
                (x"296736b5bce77ab584212116b5ad6b8420a518dce35ad9cca5"),
                (x"296736b5bce77ab584212116b5ad6b8420a518dce35ad9cca5"),
                (x"29673a528632d610ad6b5ad6b5ae105294a5295ffd2949cca5"),
                (x"29673a528632d610ad6b5ad6b5ae105294a5295ffd2949cca5"),
                (x"29673a528a52d7ded294842105294aef7b4a18dffd2949cca5"),
                (x"29673a528a52d7ded294842105294aef7b4a18dffd2949cca5"),
                (x"29673a5286377a842108e73bd31bbd421084739ce52949cca5"),
                (x"29673a5286377a842108e73bd31bbd421084739ce52949cca5"),
                (x"29673a5286377a842108e73bd31bbd421084739ce52949cca5"),
                (x"296736b5bce210f7b9ce42294a51087bdee72114a52949cca5"),
                (x"296736b5bce210f7b9ce42294a51087bdee72114a52949cca5"),
                (x"296736b5bdea10e77bdec6294e7108739def631ce35ad9cca5"),
                (x"296736b5bdea10e77bdec6294e7108739def631ce35ad9cca5"),
                (x"296736b5ad6f7a846318e71ad6b7bd42118c738d6b5ad9cca5"),
                (x"296736b5ad6f7a846318e71ad6b7bd42118c738d6b5ad9cca5"),
                (x"296736b5ad6b5b4a52946b5ad6b5ada5294a35ad6b5ad9cca5"),
                (x"296736b5ad6b5b4a52946b5ad6b5ada5294a35ad6b5ad9cca5"),
                (x"296736b5ad6b5b4a52946b5ad6b5ada5294a35ad6b5ad9cca5"),
                (x"296739ce739ce79ce7399ce739ce73ce739cce739ce739cca5"),
                (x"296739ce739ce79ce7399ce739ce73ce739cce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 12_bonus-addbomb
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739ce739ce739ce739ce739e739cce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739e739cce739cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294e739fff7b4a35ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294e739fff7b4a35ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294e739fff7b4a35ad9cca5"),
                (x"296736b5ad6f39ce739cef79ce71efef7ae710939d294ce4a5"),
                (x"296736b5ad6f39ce739cef79ce71efef7ae710939d294ce4a5"),
                (x"296736b5bce001debdef7bf9c29484ef7a4214bce35ad9cca5"),
                (x"296736b5bce001debdef7bf9c29484ef7a4214bce35ad9cca5"),
                (x"296736b5bce77ab58421842940856b10854a529ce35ad9cca5"),
                (x"296736b5bce77ab58421842940856b10854a529ce35ad9cca5"),
                (x"29673a529debde10908484294842107bdfce739ce52949cca5"),
                (x"29673a529debde10908484294842107bdfce739ce52949cca5"),
                (x"29673a529debde10908484294842107bdfce739ce52949cca5"),
                (x"29673a528f7c20b5c2107bfbda51ef739dded29ce52949cca5"),
                (x"29673a528f7c20b5c2107bfbda51ef739dded29ce52949cca5"),
                (x"29673a528f7c21083def7bdefef694a5294a529ce52949cca5"),
                (x"29673a528f7c21083def7bdefef694a5294a529ce52949cca5"),
                (x"29673a528f7bdef7bdef7bdef7bfbdef7bded29ce52949cca5"),
                (x"29673a528f7bdef7bdef7bdef7bfbdef7bded29ce52949cca5"),
                (x"29673a528633def7bdef7bdef73bbdef7b4a529ce52949cca5"),
                (x"29673a528633def7bdef7bdef73bbdef7b4a529ce52949cca5"),
                (x"29673a529ce77af7bdef7bdceef5ceef7b4a529ce52949cca5"),
                (x"29673a529ce77af7bdef7bdceef5ceef7b4a529ce52949cca5"),
                (x"29673a529ce77af7bdef7bdceef5ceef7b4a529ce52949cca5"),
                (x"296736b5bce529deb9ce73bbdef7bda5294a529ce35ad9cca5"),
                (x"296736b5bce529deb9ce73bbdef7bda5294a529ce35ad9cca5"),
                (x"296736b5bce0014a77bdef7bda5294a5294a529ce35ad9cca5"),
                (x"296736b5bce0014a77bdef7bda5294a5294a529ce35ad9cca5"),
                (x"296736b5ad6f39ce739ce739ce739ce739ce738d6b5ad9cca5"),
                (x"296736b5ad6f39ce739ce739ce739ce739ce738d6b5ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 13_bonus-power
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296736b5ad6b5ad6b5ad6b58c6b5ad6318d6b5ac635ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b58c6b5ad6318d6b5ac635ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6b58c6b5ad6318d6b5ac635ad9cca5"),
                (x"296736b5ad6b5ad6b5ad6335a6318c4210c63198c318c9cca5"),
                (x"296736b5ad6b5ad6b5ad6335a6318c4210c63198c318c9cca5"),
                (x"296736b5ad6b5ac6318c4a508631084210c621094e7399cca5"),
                (x"296736b5ad6b5ac6318c4a508631084210c621094e7399cca5"),
                (x"296736b5ad6b198c0421085084210842108421094b18c9cca5"),
                (x"296736b5ad6b198c0421085084210842108421094b18c9cca5"),
                (x"296736b5ac6630108421421080850842108421094b18c9cca5"),
                (x"296736b5ac6630108421421080850842108421094b18c9cca5"),
                (x"296736b5ac6630108421421080850842108421094b18c9cca5"),
                (x"296736b5ac65ee8477bdbdd08ef48442108421094b18c9cca5"),
                (x"296736b5ac65ee8477bdbdd08ef48442108421094b18c9cca5"),
                (x"29673631894a1084529408508a508442108421094b18c9cca5"),
                (x"29673631894a1084529408508a508442108421094b18c9cca5"),
                (x"29673631884210847bde08508ef42142108421094e7399cca5"),
                (x"29673631884210847bde08508ef42142108421094e7399cca5"),
                (x"29673631884210422108421084210842108421094b18c9cca5"),
                (x"29673631884210422108421084210842108421094b18c9cca5"),
                (x"29673ce7294a10c65294a5294a5294421084252c635ad9cca5"),
                (x"29673ce7294a10c65294a5294a5294421084252c635ad9cca5"),
                (x"29673ce7294a10c65294a5294a5294421084252c635ad9cca5"),
                (x"2967363198c21084318cce739a53184210846b4c635ad9cca5"),
                (x"2967363198c21084318cce739a53184210846b4c635ad9cca5"),
                (x"296736b5ac66b48421086318c4a5084211ad318d6b5ad9cca5"),
                (x"296736b5ac66b48421086318c4a5084211ad318d6b5ad9cca5"),
                (x"296736b5ad6b18c6210842108421296318c635ad6b5ad9cca5"),
                (x"296736b5ad6b18c6210842108421296318c635ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b18c6318c6318c6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b18c6318c6318c6b5ad6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6b18c6318c6318c6b5ad6b5ad6b5ad9cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 14_malus-inversed-commands
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"2ce739ce739ce739bdef7bdef7bdef7bdf39ce739ce739ce65"),
                (x"2ce739ce739ce739bdef7bdef7bdef7bdf39ce739ce739ce65"),
                (x"2ce739ce739ce739bdef7bdef7bdef7bdf39ce739ce739ce65"),
                (x"2ce736b5ad7bdef7ad6b5ad6b5ad6b5ad6f7bdef6b5ad9ce65"),
                (x"2ce736b5ad7bdef7ad6b5ad6b5ad6b5ad6f7bdef6b5ad9ce65"),
                (x"2ce736b5ef5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b7bdad9ce65"),
                (x"2ce736b5ef5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b7bdad9ce65"),
                (x"2ce737bd6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5adef9ce65"),
                (x"2ce737bd6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5adef9ce65"),
                (x"2ce737bd6b5ad6b5ad6b5ad6b5ad6b5ad6b5ad6b5adef9ce65"),
                (x"2ce737bd6b7bdef7ad6b5ad6b5ad6b5ad6f7bdef5adef9ce65"),
                (x"2ce737bd6b7bdef7ad6b5ad6b5ad6b5ad6f7bdef5adef9ce65"),
                (x"2bdef5adef7bdef7bdeb5ad6b5ad6b5bdef7bdef7bd6b7bde5"),
                (x"2bdef5adef7bdef7bdeb5ad6b5ad6b5bdef7bdef7bd6b7bde5"),
                (x"2bdef5adef5ad6f7bdef7bd6b5adef7bdef7ad6b7bd6b7bde5"),
                (x"2bdef5adef5ad6f7bdef7bd6b5adef7bdef7ad6b7bd6b7bde5"),
                (x"2bdef5adef5ad6f7bdef7bd6b5adef7bdef7ad6b7bd6b7bde5"),
                (x"2bdef5adef7bdef7d28f7be94a51ef7d28f7bdef7bd6b7bde5"),
                (x"2bdef5adef7bdef7d28f7be94a51ef7d28f7bdef7bd6b7bde5"),
                (x"2bdef5ad6b7bdef7d28b5ae94a516b5d28f7bdef5ad6b7bde5"),
                (x"2bdef5ad6b7bdef7d28b5ae94a516b5d28f7bdef5ad6b7bde5"),
                (x"2bdef5ad6b5ad6b5d294a5294a5294a528b5ad6b5ad6b7bde5"),
                (x"2bdef5ad6b5ad6b5d294a5294a5294a528b5ad6b5ad6b7bde5"),
                (x"2bdef5ad6b5ad6b5d294a5294a5294a528b5ad6b5ad6b7bde5"),
                (x"2ce737bd6b5ad6b5ad6b5ae94a516b5ad6b5ad6b5adef9ce65"),
                (x"2ce737bd6b5ad6b5ad6b5ae94a516b5ad6b5ad6b5adef9ce65"),
                (x"2ce736b5ef7bdeb5ad6b5ae94a516b5ad6b5bdef7bdad9ce65"),
                (x"2ce736b5ef7bdeb5ad6b5ae94a516b5ad6b5bdef7bdad9ce65"),
                (x"2ce736b5ad7bdeb5d294a5294a5294a528b5bdef6b5ad9ce65"),
                (x"2ce736b5ad7bdeb5d294a5294a5294a528b5bdef6b5ad9ce65"),
                (x"2ce736b5ad7bdeb5d294a5294a5294a528b5bdef6b5ad9ce65"),
                (x"2ce736b5ad7bdeb5d28b5adef7bd6b5d28b5bdef6b5ad9ce65"),
                (x"2ce736b5ad7bdeb5d28b5adef7bd6b5d28b5bdef6b5ad9ce65"),
                (x"2ce736b5ad7bdf4a528f7bdef7bdef7d294a3def6b5ad9ce65"),
                (x"2ce736b5ad7bdf4a528f7bdef7bdef7d294a3def6b5ad9ce65"),
                (x"2ce739ce739ce739ce739ce739ce739ce739ce739ce739ce65"),
                (x"2ce739ce739ce739ce739ce739ce739ce739ce739ce739ce65"),
                (x"2ce739ce739ce739ce739ce739ce739ce739ce739ce739ce65"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 15_malus-disable-bombs
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce79ce7339ce73ce694a53399ce739e739cce739cca5"),
                (x"296739ce79ce7339ce73ce694a53399ce739e739cce739cca5"),
                (x"29739a5294a529ded294a510818e94a529ded294a5294ce4a5"),
                (x"29739a5294a529ded294a510818e94a529ded294a5294ce4a5"),
                (x"29739a5294a529ded294a510818e94a529ded294a5294ce4a5"),
                (x"29739a528840c7ce1ce739c21423bd00014a0c6845294ce4a5"),
                (x"29739a528840c7ce1ce739c21423bd00014a0c6845294ce4a5"),
                (x"29673a528319cf0877bd18c2142063a5280077a31d2949cca5"),
                (x"29673a528319cf0877bd18c2142063a5280077a31d2949cca5"),
                (x"29673e739ce2d6b5d29418d0842063a529ded29ce77bd9cca5"),
                (x"29673e739ce2d6b5d29418d0842063a529ded29ce77bd9cca5"),
                (x"29673a529ffad610c21018d0842063a529ded280052949cca5"),
                (x"29673a529ffad610c21018d0842063a529ded280052949cca5"),
                (x"29673a529ffad610c21018d0842063a529ded280052949cca5"),
                (x"29673a529082d61084217be94a53de739dded29ce52949cca5"),
                (x"29673a529082d61084217be94a53de739dded29ce52949cca5"),
                (x"29673a529083def7ad6b5ae10841efef7bce5280052949cca5"),
                (x"29673a529083def7ad6b5ae10841efef7bce5280052949cca5"),
                (x"29673a528e70c74a3def842107bdcea5294a0c74a52949cca5"),
                (x"29673a528e70c74a3def842107bdcea5294a0c74a52949cca5"),
                (x"29739a528318428452947bdef73b9ca5288404231d294ce4a5"),
                (x"29739a528318428452947bdef73b9ca5288404231d294ce4a5"),
                (x"29739a52810842845294ef7bdef694a5288404210d294ce4a5"),
                (x"29739a52810842845294ef7bdef694a5288404210d294ce4a5"),
                (x"29739a52810842845294ef7bdef694a5288404210d294ce4a5"),
                (x"29739a528840c631d294a5294a5294a528318c6845294ce4a5"),
                (x"29739a528840c631d294a5294a5294a528318c6845294ce4a5"),
                (x"296736b5bce0014a5294a5294a5294a5294a001ce35ad9cca5"),
                (x"296736b5bce0014a5294a5294a5294a5294a001ce35ad9cca5"),
                (x"296736b5ad6f39ce739ce739ce739ce739ce738d6b5ad9cca5"),
                (x"296736b5ad6f39ce739ce739ce739ce739ce738d6b5ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"296736b5ad6b5ad6d294a5294a5294a528d6b5ad6b5ad9cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),

                -- 16_malus-remove-power
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739b5ad6b5ad6b58c6b5ad6318c64e739ce739cca5"),
                (x"296739ce739b5ad6b5ad6b58c6b5ad6318c64e739ce739cca5"),
                (x"296739ce739b5ad6b5ad6b58c6b5ad6318c64e739ce739cca5"),
                (x"296739ce739ce6d6b5ad6335a6318cc63139ce739ce739cca5"),
                (x"296739ce739ce6d6b5ad6335a6318cc63139ce739ce739cca5"),
                (x"296739ce739ce739b18c4a508631299ce739ce739e7399cca5"),
                (x"296739ce739ce739b18c4a508631299ce739ce739e7399cca5"),
                (x"29673f7bd39ce739ce73bdd084a6739ce739ce694b18c9cca5"),
                (x"29673f7bd39ce739ce73bdd084a6739ce739ce694b18c9cca5"),
                (x"296736b5b9cce739ce739cd299ce739ce739a1094b18c9cca5"),
                (x"296736b5b9cce739ce739cd299ce739ce739a1094b18c9cca5"),
                (x"296736b5b9cce739ce739cd299ce739ce739a1094b18c9cca5"),
                (x"296736b5ac656b39ce739ce739ce739ce68421094b18c9cca5"),
                (x"296736b5ac656b39ce739ce739ce739ce68421094b18c9cca5"),
                (x"29673631894a1094ce739ce739ce7342108421094b18c9cca5"),
                (x"29673631894a1094ce739ce739ce7342108421094b18c9cca5"),
                (x"29673631884210844e739ce739ce734a528421094e7399cca5"),
                (x"29673631884210844e739ce739ce734a528421094e7399cca5"),
                (x"2967363188421139ce739ce739ce739ce694a1094b18c9cca5"),
                (x"2967363188421139ce739ce739ce739ce694a1094b18c9cca5"),
                (x"29673ce7294ce739ce739cd8c9ce739ce739eb4c635ad9cca5"),
                (x"29673ce7294ce739ce739cd8c9ce739ce739eb4c635ad9cca5"),
                (x"29673ce7294ce739ce739cd8c9ce739ce739eb4c635ad9cca5"),
                (x"29673631939ce739ce739cf39a52739ce739ce79cb5ad9cca5"),
                (x"29673631939ce739ce739cf39a52739ce739ce79cb5ad9cca5"),
                (x"296739ce739ce739a5296318c4a5089ce739ce739b18c9cca5"),
                (x"296739ce739ce739a5296318c4a5089ce739ce739b18c9cca5"),
                (x"296739ce739ce79ca1084210842129631939ce739ce739cca5"),
                (x"296739ce739ce79ca1084210842129631939ce739ce739cca5"),
                (x"296739ce739b18d6b18c6318c6318c6b5ad6ce739ce739cca5"),
                (x"296739ce739b18d6b18c6318c6318c6b5ad6ce739ce739cca5"),
                (x"296739ce739b18d6b18c6318c6318c6b5ad6ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"296739ce739ce739ce739ce739ce739ce739ce739ce739cca5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5"),
                (x"294a5294a5294a5294a5294a5294a5294a5294a5294a5294a5")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 1679 := 0;
    signal out_color_reg : std_logic_vector(199 downto 0) := (others => '0');
begin
    process(in_sprite_id, in_sprite_row, in_sprite_col, in_sprite_state, in_sprite_direction)
    begin
        real_row <= 0;
        case in_sprite_id is
            when 0 => real_row <= in_sprite_row;
            when 1 => real_row <= 40 + in_sprite_row;
            when 2 => real_row <= 80 + in_sprite_row;
            when 3 => real_row <= 120 + in_sprite_row;
            when 4 =>
                case in_sprite_state is
                    when 0 => real_row <= 160 + in_sprite_row;
                    when others => null;
                end case;
            when 5 =>
                case in_sprite_state is
                    when 0 => real_row <= 200 + in_sprite_row;
                    when 1 => real_row <= 240 + in_sprite_row;
                    when 2 => real_row <= 280 + in_sprite_row;
                    when 3 => real_row <= 320 + in_sprite_row;
                    when others => null;
                end case;
            when 6 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 360 + in_sprite_row;
                            when D_LEFT => real_row <= 400 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 440 + in_sprite_row;
                            when D_LEFT => real_row <= 480 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 520 + in_sprite_row;
                            when D_LEFT => real_row <= 560 + in_sprite_row;
                            when others => null;
                        end case;
                    when 3 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 600 + in_sprite_row;
                            when D_LEFT => real_row <= 640 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 7 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 680 + in_sprite_row;
                            when D_LEFT => real_row <= 720 + in_sprite_row;
                            when D_DOWN => real_row <= 760 + in_sprite_row;
                            when D_RIGHT => real_row <= 800 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 840 + in_sprite_row;
                            when D_LEFT => real_row <= 880 + in_sprite_row;
                            when D_DOWN => real_row <= 920 + in_sprite_row;
                            when D_RIGHT => real_row <= 960 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1000 + in_sprite_row;
                            when D_LEFT => real_row <= 1040 + in_sprite_row;
                            when D_DOWN => real_row <= 1080 + in_sprite_row;
                            when D_RIGHT => real_row <= 1120 + in_sprite_row;
                            when others => null;
                        end case;
                    when 3 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1160 + in_sprite_row;
                            when D_LEFT => real_row <= 1200 + in_sprite_row;
                            when D_DOWN => real_row <= 1240 + in_sprite_row;
                            when D_RIGHT => real_row <= 1280 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 8 => real_row <= 1320 + in_sprite_row;
            when 9 => real_row <= 1360 + in_sprite_row;
            when 10 => real_row <= 1400 + in_sprite_row;
            when 11 => real_row <= 1440 + in_sprite_row;
            when 12 => real_row <= 1480 + in_sprite_row;
            when 13 => real_row <= 1520 + in_sprite_row;
            when 14 => real_row <= 1560 + in_sprite_row;
            when 15 => real_row <= 1600 + in_sprite_row;
            when 16 => real_row <= 1640 + in_sprite_row;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= rom(real_row);
        end if;
    end process;
    out_color <= out_color_reg(((in_sprite_col + 1) * 5) - 1 downto (in_sprite_col * 5));
end behavioral;
