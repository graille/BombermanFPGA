library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_nb : in integer range 0 to 52;
        in_sprite_row : in integer range 0 to 66;
        in_sprite_col : in integer range 0 to 39;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end sprite_rom;

architecture behavioural of sprite_rom is
    subtype word_t is std_logic_vector(39 downto 0);
    type memory_t is array(2515 downto 0) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- block.bmp
                ("00110001100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000111001110011100011000110001100011000110001100011000110001100011"),
                ("00110001100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000111001110011100011000110001100011000110001100011000110001100011"),
                ("00111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001100011000111001110011100111001110011100111001110011100111001110011100111"),
                ("00111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001100011000111001110011100111001110011100111001110011100111001110011100111"),
                ("00111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001100011000111001110011100111001110011100111001110011100111001110011100111"),
                ("00110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("00110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("00101001010010100101001010010100101001100011000110001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100001100011000110010100101"),
                ("00101001010010100101001010010100101001100011000110001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100001100011000110010100101"),
                ("00101001010010100101001010010100101001100011000110001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100001100011000110010100101"),
                ("00101001010010100101001010010100101001100011000110001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110001100011000110010100101"),
                ("00101001010010100101001010010100101001100011000110001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110001100011000110010100101"),
                ("00011000110001100011000110001100011001110011100111001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110001100011000110001100011"),
                ("00011000110001100011000110001100011001110011100111001010010100101001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110001100011000110001100011"),
                ("00011000110001100011000110001100011001100011000110001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100111001110001100011000110001100011"),
                ("00011000110001100011000110001100011001100011000110001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100111001110001100011000110001100011"),
                ("00011000110001100011000110001100011001100011000110001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100111001110001100011000110001100011"),
                ("00111001110011000110001100011000110001100011000110001100011000110001110011100110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000111001110011100111001110011100111"),
                ("00111001110011000110001100011000110001100011000110001100011000110001110011100110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000111001110011100111001110011100111"),
                ("00100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000100001000010000100001000010000100"),
                ("00100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000100001000010000100001000010000100"),
                ("00100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000100001000010000100001000010000100"),
                ("00100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000100001000010000100001000010000100"),
                ("00100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000100001000010000100001000010000100"),
                ("00100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000100001000010000100001000010000100"),
                ("00101001010010100101001010010100101001010010100101001010010100101001010010100111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000101001010010100101001010010100101"),
                ("00101001010010100101001010010100101001010010100101001010010100101001010010100111001110011100011000110001100011000110001100011000110001100011000110001100110001100011000101001010010100101001010010100101"),
                ("00111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000111001110011100111001110011100111"),
                ("00111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000111001110011100111001110011100111"),
                ("00111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000111001110011100111001110011100111"),
                ("00110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("00110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),

                -- bomb_1_0.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100100001001110111101111011110111101001000010000100000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100100001001110111101111011110111101001000010000100000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000110001100011000011000110001100011000110001100011000110001100011001100011000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000110001100011000011000110001100011000110001100011000110001100011001100011000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100110001100000000000000001111111111111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111111111011110111100000000000000000011000110001100011000110001100011000111001110011100111001110011100111001110011100111001100011000110001100011000110001100000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011000110001100011000110001100011000111001110011100111001110011100111001110011100111001100011000110001100011000110001100000000000000001111011110111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- bomb_1_1.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100110100001000010001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100110100001000010001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000001001110011100111001110011000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000001001110011100111001110011000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100100001001110111101111011110111101001000010000100000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100100001001110111101111011110111101001000010000100000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000110001100011000011000110001100011000110001100011000110001100011001100011000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000110001100011000011000110001100011000110001100011000110001100011001100011000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100110001100000000000000001111111111111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111111111011110111100000000000000000011000110001100011000110001100011000111001110011100111001110011100111001110011100111001100011000110001100011000110001100000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011000110001100011000110001100011000111001110011100111001110011100111001110011100111001100011000110001100011000110001100000000000000001111011110111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- bomb_1_2.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111110011100111100011000110001100011000100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001111000110001100011000110000100001000110001100011000100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001111000110001100011000110000100001000110001100011000100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001111000110001100011000110000100001000110001100011000100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001111000110000100001000010000100001000110001100011000100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001111000110000100001000010000100001000110001100011000100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001110011100111100011000110001100011000100111001110011100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001110011100111100011000110001100011000100111001110011100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111110011100111001110011100111100011000110001100011000100111001110011100111001111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111010011100111001110011100111001110011100111001110011111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111010011100111001110011100111001110011100111001110011111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111000000000000000000100001001110111101111011110111101001000010000100000000000011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100100001001110111101111011110111101001000010000100000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100100001001110111101111011110111101001000010000100000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111000000000000011000110001100011000110010000100001000010000100000110001100011000110001100000000000000011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000110001100011000011000110001100011000110001100011000110001100011001100011000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000110001100011000011000110001100011000110001100011000110001100011001100011000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100110001100000000000000001111111111111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011100111001110011100111001110011100111001111000010000100001000010000001110011100111001110011100111001110011100111001110000000000000001111011110111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111110000000000000000011000110001100011000110001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001100000000000111111111111111"),
                ("11111111111111011110111100000000000000000011000110001100011000110001100011000111001110011100111001110011100111001110011100111001100011000110001100011000110001100000000000000001111011110111111111111111"),
                ("11111111111111011110111100000000000000000011000110001100011000110001100011000111001110011100111001110011100111001110011100111001100011000110001100011000110001100000000000000001111011110111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111110000000000000000011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100000000000000001111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011110111100000000000001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000000000001111011110111101111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011110000000000000000000000000000110001100011000110001100011000110001100011000110000000000000000000000000011110111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111110111101111000000000000000000000000000000000000000000000000000111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- bonus_bomb.bmp
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010010100101001010001101011011010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010010100101001010001101011011010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010010100101001010001101011011010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010010100101001010001110011100111001110101001010010100011110111101110011100111010100101000000100001000011001110011101001010010011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010010100101001010001110011100111001110101001010010100011110111101110011100111010100101000000100001000011001110011101001010010011100111001101011"),
                ("10011100110110101101011011010010100101001010010100011100111001111011110111101111011111010010100100001000010000000010000110100101001010000001000011000010000100001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100011100111001111011110111101111011111010010100100001000010000000010000110100101001010000001000011000010000100001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100011100111001111011110111101111011111010010100100001000010000000010000110100101001010000001000011000010000100001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100011100111001110100001000000001000010000110000100001010010100000010000100001000010000110100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100011100111001110100001000000001000010000110000100001010010100000010000100001000010000110100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100111010010100101001010010100011110111101111000010000100001000010000110000100001010010100100001000010000100001000001111011110111101110011100111001110011101010010100101001010010011100111001101011"),
                ("10011100111010010100101001010010100011110111101111000010000100001000010000110000100001010010100100001000010000100001000001111011110111101110011100111001110011101010010100101001010010011100111001101011"),
                ("10011100111010010100101001010010100011110111101111000010000100001000010000110000100001010010100100001000010000100001000001111011110111101110011100111001110011101010010100101001010010011100111001101011"),
                ("10011100111010010100101000111001110100001000010000010110101110000100001000001111011110111001110101001010010100011110111101110011100111001110011101010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111001110100001000010000010110101110000100001000001111011110111001110101001010010100011110111101110011100111001110011101010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111101111011110111101111100001000001111011110111101111011110111101111011100111001110101001010010100101001010010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111101111011110111101111100001000001111011110111101111011110111101111011100111001110101001010010100101001010010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111101111011110111101111011110111101111011110111101111011110111101111011110111101111011100111001110011100111001110011101010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111101111011110111101111011110111101111011110111101111011110111101111011110111101111011100111001110011100111001110011101010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111101111011110111101111011110111101111011110111101111011110111101111011110111101111011100111001110011100111001110011101010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111001110011110111101111011110111101111011110111101111011110111101111011100111001110011100111001110011100111010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101000111001110011110111101111011110111101111011110111101111011110111101111011100111001110011100111001110011100111010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101001010010100011100111001110011110111101111011110111101111011110111001110011100111001110011100111001110011100111010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101001010010100011100111001110011110111101111011110111101111011110111001110011100111001110011100111001110011100111010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100111010010100101001010010100011100111001110011110111101111011110111101111011110111001110011100111001110011100111001110011100111010100101001010010100101001010010100101001010010011100111001101011"),
                ("10011100110110101101011011010010100101001010010100011100111001110011100111001110011100111001110011100111001110011100111010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100011100111001110011100111001110011100111001110011100111001110011100111010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100101001010001110011100111001110011100111001110101001010010100101001010010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100101001010001110011100111001110011100111001110101001010010100101001010010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100101001010001110011100111001110011100111001110101001010010100101001010010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010010100101001010001101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010010100101001010001101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("01011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011"),

                -- bonus_life.bmp
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100101001010010100101001010010100101000110101101011010110101101101001010010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100101001010010100101001010010100101000110101101011010110101101101001010010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100101001010010100101001010010100101001010010100101000110101101011010110101101101001010010100101001010010100101001010010100101001010010100011010110110011100111001101011"),
                ("10011100111010010100101000110001100100111001110011010010100110011100111001101100011001010010100101001010010100011000110010011100111001110011100111001110011100110110001100101001010010011100111001101011"),
                ("10011100111010010100101000110001100100111001110011010010100110011100111001101100011001010010100101001010010100011000110010011100111001110011100111001110011100110110001100101001010010011100111001101011"),
                ("10100101000110001100011001001110011010000100001000000010000101001010010100110011100110110001100011000110001100100111001110011100111001101001010011001110011100111001110011011000110010100101001010001011"),
                ("10100101000110001100011001001110011010000100001000000010000101001010010100110011100110110001100011000110001100100111001110011100111001101001010011001110011100111001110011011000110010100101001010001011"),
                ("10100101000110001100011001001110011010000100001000000010000101001010010100110011100110110001100011000110001100100111001110011100111001101001010011001110011100111001110011011000110010100101001010001011"),
                ("10100101000110001100011000100101001000010000100001010000100001001010010100110100101001001110011100111001110011101001010001001010010100101001010010100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100101001000010000100001010000100001001010010100110100101001001110011100111001110011101001010001001010010100101001010010100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100001000000010000100001010000100001001010010100110100101000100101001010010100101001101001010001001010010100101000010000100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100001000000010000100001010000100001001010010100110100101000100101001010010100101001101001010001001010010100101000010000100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100001000000010000100001010000100001001010010100110100101000100101001010010100101001101001010001001010010100101000010000100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100001000010000100001000010000100001000010000100010100101000100101001010010100101001101001010001000010000100001000010000100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100001000010000100001000010000100001000010000100010100101000100101001010010100101001101001010001000010000100001000010000100101001010011001110011011000110010100101001010001011"),
                ("10100101000110001100011000100101001010000100001000010000100001001010010100110100101000100101001010010100101001101001010001000010000100001001010011001110011100111001110011011000110010100101001010001011"),
                ("10100101000110001100011000100101001010000100001000010000100001001010010100110100101000100101001010010100101001101001010001000010000100001001010011001110011100111001110011011000110010100101001010001011"),
                ("10011100111010010100101001001110011010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010011001110011100111001110011101001010010011100111001101011"),
                ("10011100111010010100101001001110011010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010011001110011100111001110011101001010010011100111001101011"),
                ("10011100111010010100101001001110011010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010011001110011100111001110011101001010010011100111001101011"),
                ("10011100111010010100101000110001100010010100101001010010100110100101001010010011100110100101001010010100101001100111001110100101001010010011100111001110011100110110001100101001010010011100111001101011"),
                ("10011100111010010100101000110001100010010100101001010010100110100101001010010011100110100101001010010100101001100111001110100101001010010011100111001110011100110110001100101001010010011100111001101011"),
                ("10011100110110101101011011010010100011000110001100010010100110011100111001110100101001010010100101001010010100101001010010011100111001110011100110110001100011001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100011000110001100010010100110011100111001110100101001010010100101001010010100101001010010011100111001110011100110110001100011001010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100011000110001100010010100110011100111001110100101001010010100101001010010100101001010010011100111001110011100110110001100011001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100011000110010011100111001101001010010100101001010010100101001100111001110011100111001101100011001010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100011000110010011100111001101001010010100101001010010100101001100111001110011100111001101100011001010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010010011100110100101001100111001110011100111001110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010010011100110100101001100111001110011100111001110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010010011100110100101001100111001110011100111001110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101001001110011100111001110011101001010001101011010110101101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101001001110011100111001110011101001010001101011010110101101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110101101011011010010100101001010010100011010110101101011010110101101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110101101011011010010100101001010010100011010110101101011010110101101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("01011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011"),

                -- bonus_power.bmp
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110101101011011010010100011010110101101011010110110100101001010001101011010110101101011011010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110101101011011010010100011010110101101011010110110100101001010001101011010110101101011011010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110101101011011010010100011010110101101011010110110100101001010001101011010110101101011011010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000100101001101001010010100101001010001001010010100110100101001010010100101001001110011101001010010011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000100101001101001010010100101001010001001010010100110100101001010010100101001001110011101001010010011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010001001010010100001000101001010010100010010100101000010000100010100101000100101001010010100101001101001010010011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010001001010010100001000101001010010100010010100101000010000100010100101000100101001010010100101001101001010010011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010001001010010100001000101001010010100010010100101000010000100010100101000100101001010010100101001101001010010011100111001101011"),
                ("10011100110110101101011010110101101101001010010100010010100101000010000100000001000010100001000010010100101001000010000101000010000100001001010010100001000010000100101001101001010010011100111001101011"),
                ("10011100110110101101011010110101101101001010010100010010100101000010000100000001000010100001000010010100101001000010000101000010000100001001010010100001000010000100101001101001010010011100111001101011"),
                ("10011100110110101101011011010010100010010100101001010000100000001000010000101000010000100001000010000100001000000010000101000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100110110101101011011010010100010010100101001010000100000001000010000101000010000100001000010000100001000000010000101000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100110110101101011011010010100010010100101001010000100000001000010000101000010000100001000010000100001000000010000101000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100110110101101011011010010100010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100110110101101011011010010100010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100111010010100101000100101001010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100111010010100101000100101001010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100111010010100101000100001000010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100111010010100101000100001000010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100111010010100101000100001000010000100001000000010000110100101001010001000010000100001000101001010010100010000100001000010000100001000010000100001000010000100101001101001010010011100111001101011"),
                ("10011100111010010100101000100001000010000100001000010000100000001000010000101000010000100001000010000100001000010000100001000010000100001000010000100001000010001001110011101001010010011100111001101011"),
                ("10011100111010010100101000100001000010000100001000010000100000001000010000101000010000100001000010000100001000010000100001000010000100001000010000100001000010001001110011101001010010011100111001101011"),
                ("10011100111010010100101000100101001010000100001000101001010010100101001010010100101001010010100101001010010100101001010001000010000100001000010000100101001010011010010100011010110110011100111001101011"),
                ("10011100111010010100101000100101001010000100001000101001010010100101001010010100101001010010100101001010010100101001010001000010000100001000010000100101001010011010010100011010110110011100111001101011"),
                ("10011100111010010100101000100101001010000100001000101001010010100101001010010100101001010010100101001010010100101001010001000010000100001000010000100101001010011010010100011010110110011100111001101011"),
                ("10011100111010010100101001001110011010000100001000010000100010100101001010010011100111001110011101001010010100010010100101000010000100001001010011001110011100111010010100011010110110011100111001101011"),
                ("10011100111010010100101001001110011010000100001000010000100010100101001010010011100111001110011101001010010100010010100101000010000100001001010011001110011100111010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100100111001110011010010100101000010000100010100101001010010100010010100101001010000100001001010010100110011100111010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011011010010100100111001110011010010100101000010000100010100101001010010100010010100101001010000100001001010010100110011100111010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011011010010100100111001110011010010100101000010000100010100101001010010100010010100101001010000100001001010010100110011100111010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010001001010010100101000010000100001000010000100001000100111001110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010001001010010100101000010000100001000010000100001000100111001110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010001101011010110101101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010010100101001010010100101001010010100101001010001101011010110101101011010110101101011010110101101011010110110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("01011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011"),

                -- bonus_speed.bmp
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000110001100011000110001100011000110001100011000110001100011000110001100011001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000110001100011000110001100011000110001100011000110001100011000110001100011001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000110001100011000110001100011000110001100011000110001100011000110001100011001010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101001000010000000010000100001010110101110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101001000010000000010000100001010110101110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010001000010000100001000010010100101001100111001110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010001000010000100001000010010100101001100111001110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010001000010000100001000010010100101001100111001110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000101001010010100101001010010100101010000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110101101011010110110100101000101001010010100101001010010100101010000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010001000010000100001000010010100101001100111001110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010001000010000100001000010010100101001100111001110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101011010110110100101001010001000010000100001000010010100101001100111001110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010010100101001010010100101000101001010010100101001010010100101010000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100101001010010100101001010010100101000101001010010100101001010010100101010000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100011100111001110010110101100001000010000100001000010101101011010110101101011010110101110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100011100111001110010110101100001000010000100001000010101101011010110101101011010110101110000100001000001010010100111001110011101010010100011010110110011100111001101011"),
                ("10011100111010010100101000111001110010110101101011000010000101011010110101101011010110101101011010110101101011100001000001010010100101001010010100101001010010100111001110101001010010011100111001101011"),
                ("10011100111010010100101000111001110010110101101011000010000101011010110101101011010110101101011010110101101011100001000001010010100101001010010100101001010010100111001110101001010010011100111001101011"),
                ("10011100111010010100101000111001110010110101101011000010000101011010110101101011010110101101011010110101101011100001000001010010100101001010010100101001010010100111001110101001010010011100111001101011"),
                ("10011100111010010100101000101001010010110101101011101001010010100101001010010000100001000010000010100101001010010100101010100101001010010100101000111001110011100111001110101001010010011100111001101011"),
                ("10011100111010010100101000101001010010110101101011101001010010100101001010010000100001000010000010100101001010010100101010100101001010010100101000111001110011100111001110101001010010011100111001101011"),
                ("10011100111010010100101000111001110101001010010100010000100001000010000100010100101000111001110011100111001110101001010001000010000100001000010001010010100101000111001110101001010010011100111001101011"),
                ("10011100111010010100101000111001110101001010010100010000100001000010000100010100101000111001110011100111001110101001010001000010000100001000010001010010100101000111001110101001010010011100111001101011"),
                ("10011100111010010100101000111001110101001010010100010000100001000010000100010100101000111001110011100111001110101001010001000010000100001000010001010010100101000111001110101001010010011100111001101011"),
                ("10011100110110101101011011010010100010000100001000011110111101110011100111001000010001010010100101001010010100010000100001111011110111101110011100100001000010001010010100101001010010011100111001101011"),
                ("10011100110110101101011011010010100010000100001000011110111101110011100111001000010001010010100101001010010100010000100001111011110111101110011100100001000010001010010100101001010010011100111001101011"),
                ("10011100110110101101011011010010100010000100001000011100111001110011100111001001010011010010100101001010010100010000100001110011100111001110011100100101001010011010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100010000100001000011100111001110011100111001001010011010010100101001010010100010000100001110011100111001110011100100101001010011010010100011010110110011100111001101011"),
                ("10011100110110101101011011010010100010000100001000011100111001110011100111001001010011010010100101001010010100010000100001110011100111001110011100100101001010011010010100011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100010000100001001010010100110100101000110101101011010110101101101001010001000010000100001001010011010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101101001010010100010000100001001010010100110100101000110101101011010110101101101001010001000010000100001001010011010010100101000110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010001101011010110101101011010110101101011010110110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100110110101101011010110101101011010110101101101001010010100101001010001101011010110101101011010110101101011010110110100101001010010100101000110101101011010110101101011010110110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("10011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001101011"),
                ("01011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011"),

                -- character_D_0.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000001000010010000100010100101011100111001110001000010000100001000111001110011100010100101000100001000000100001111001110011100111001111111111111111111111111"),
                ("11111111111111111111111001101011010110101101011010110101110011100010100101001010010100101001010010100101001010010100101001010010100101011100111001101011010110101101011010110101110011111111111111111111"),
                ("11111111111111111111111001101011010110101101011010110101110011100010100101001010010100101001010010100101001010010100101001010010100101011100111001101011010110101101011010110101110011111111111111111111"),
                ("11111111111111111111111001101011010100111001110011100111110011100001000010001010010100101001010010100101001010010100101001010001000010011100111001001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111001101011010100111001110011100111110011100001000010001010010100101001010010100101001010010100101001010001000010011100111001001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111110011100001000010000100111001110011100111001110011100111001110000100001000010011100111001001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111110011100001000010000100111001110011100111001110011100111001110000100001000010011100111001001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111111110011100111001110011100111001110011100001000010000100111001110011111111111111111111111001110000100001000010011100111001110011100111001110011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011100111001110011100001000010000100111001110011111111111111111111111001110000100001000010011100111001110011100111001110011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011111111111111111111111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010100111001110011111001110011111111111111111111111001110010011100111001111010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010100111001110011111001110011111111111111111111111001110010011100111001111010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011111001110011111111111111111111111001110010011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011111001110011111111111111111111111001110010011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011100111001111010111001110011111111111111111111111001110011010100111001110011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011100111001111010111001110011111111111111111111111001110011010100111001110011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010110101101011100111111111111111111111111111111111111111111100110101101011010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010110101101011100111111111111111111111111111111111111111111100110101101011010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_D_1.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010001010010100100001000010000100001010010101010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010001010010100100001000010000100001010010101010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100010100101001010010100101001010010100101001010010100101001010010100101011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100010100101001010010100101001010010100101001010010100101001010010100101011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101101011010110101101011100111001110001000010000100001000111001110011100010100101011100111001101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101101011010110101101011100111001110001000010000100001000111001110011100010100101011100111001101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011110101101001010010100101001010010100101001010010100101001010111001110010011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011110101101001010010100101001010010100101001010010100101001010111001110010011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001100100010100101001010010100101001010001000010000100111001110010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001100100010100101001010010100101001010001000010000100111001110010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100001000010000100111001110011100111001110011100001000010000100111001110011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100001000010000100111001110011100111001110011100001000010000100111001110011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100001000010011100111000010000100100111001111010100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001100100001000010011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001100100001000010011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010100111001110011110101101011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010100111001110011110101101011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011110101101011010110101101010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011110101101011010110101101010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_D_2.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010110101101011010100111001101010010100101001010010100101001010010100101011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010110101101011010100111001101010010100101001010010100101001010010100101011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011110101101010011100111001101010010100101001010010100101001010111001110011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011110101101010011100111001101010010100101001010010100101001010111001110011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001101000010000100001000111001110011100010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001101000010000100001000111001110011100010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100001000010011100010100101001010010100101001010100111001110011110101101010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011100111001001110011100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011100111001001110011100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010100111001100100111001110011100111001001110011110101101011010110101101011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010100111001100100111001110011100111001001110011110101101011010110101101011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_D_4.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100010100101001010010100101001010010100101001010100111001111010110101101011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100010100101001010010100101001010010100101001010100111001111010110101101011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100111001110001010010100101001010010100101001010100111001110011110101101010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100111001110001010010100101001010010100101001010100111001110011110101101010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101011100111001110001000010000100001000100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101011100111001110001000010000100001000100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011110101101010011100111001101010010100101001010010100101011100001000010000100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001110011100111110011100111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001110011100111110011100111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010110101101011010110101101010011100111110011100111001110000100100111001111010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010110101101011010110101101010011100111110011100111001110000100100111001111010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001110011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001110011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_D_5.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001111010110101101011010100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000110111101111011110111101111011110111101111011110111000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000011011110111101111011110111101111011110111101111011110111101111011110111101111011110111101110000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011100001101111011110111101111011110111101111011100001101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000110111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010010111101111011110111101111011111100101111011110111101111011110111101111011111100101111011110111101111011110111001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110001001010011011110111101111011111100101111011110111101111011110111101111011111100101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000100101001010010100101001101111011110111101111011110111101111011101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010101001010010100101001010010100101001010010100101001001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010001010010100100001000010000100001010010101010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010001010010100100001000010000100001010010101010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100010100101001010010100101001010010100101001010010100101001010010100101000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100010100101001010010100101001010010100101001010010100101001010010100101000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101110011100010100101011100111001110001000010000100001000111001110011100110101101011010110101101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101110011100010100101011100111001110001000010000100001000111001110011100110101101011010110101101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011111001110001010010100101001010010100101001010010100101001010110101101010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011111001110001010010100101001010010100101001010010100101001010110101101010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011111001110000100001000010001010010100101001010010100101000100100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011111001110000100001000010001010010100101001010010100101000100100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100111001110000100001000010011100111001110011100111001110000100001000010011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100111001110000100001000010011100111001110011100111001110000100001000010011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001111010100111001100100001001110011100001000010000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100001000010000100100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100001000010000100100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100110101101010011100111001111010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100110101101010011100111001111010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011110101101011010110101101010011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011110101101011010110101101010011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_R_0.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011110101101011010110101001110011111001110011111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011110101101011010110101001110011111001110011111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110000100001001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110000100001001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000100001000010000100001101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000100001000010000100001101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011110111101111011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011110111101111011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011100001000011011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011100001000011011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000011011110111101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000011011110111101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001010010100101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110001010001000010000001000010101001010010100101001010010000100011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110001010001000010000001000010101001010010100101001010010000100011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101011100001000010000001000011110011100111001110011100010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110001010110101101011010110101101011010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110001010110101101011010110101101011010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111101011010010100101011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111101011010010100101011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000100001000010000100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000100001000010000100100111001111010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000100001000010000100100111001111010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100100111001110011100111001110011100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100110101101010011100111001110011100111001110011110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111100110101101010011100111001110011100111001110011110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011010110101101011010110101101011010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011010110101101011010110101101011010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_R_1.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011110101101011010110101001110011111001110011111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011110101101011010110101001110011111001110011111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110000100001001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110000100001001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000100001000010000100001101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000100001000010000100001101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011110111101111011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011110111101111011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011100001000011011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011100001000011011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000011011110111101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000011011110111101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001010010100101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001000010000001000010101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110000100000010000101010010100101001010010100101001010010000100011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110000100000010000101010010100101001010010100101001010010000100011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010110101101011010000010000111100111001110011100111001110011100010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001111010010100101001010010100101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001111010010100101001010010100101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000101001011110011100111001110011100111001110000100001000010000100001000010011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000101001011110011100111001110011100111001110000100001000010000100001000010011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110010100101001010010111100111001110000100001000010000100001000010011100111111111111100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110010100101001010010111100111001110000100001000010000100001000010011100111111111111100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111001110011100111001110011111001110011100111000010000100001000010000100111001110011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111001110011100111001110011100111001111100111000010000100001000010000100100111001110011100111001110011100111001111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111001110011100111001110011100111001111100111000010000100001000010000100100111001110011100111001110011100111001111100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001111100111001110011100001000010010011100111001110011100111001110011110101101011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001111100111001110011100001000010010011100111001110011100111001110011110101101011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100100111001110011111001110011111111111110011100100111001110011100111001111010110101101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100100111001110011111001110011111111111110011100100111001110011100111001111010110101101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100110101101011010110101101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100110101101011010110101101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_R_2.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011110101101011010110101001110011111001110011111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011110101101011010110101001110011111001110011111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110000100001001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100110000100001001000010000001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000100001000010000100001101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000100001000010000100001101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011110111101111011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011110111101111011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011100001000011011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011100001000011011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000011011110111101111011110111101111011111100111001011110111111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000011011110111101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000011011110111101111011110111101111011110111101110100101001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001010010100101001010010100101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101000001000010000100100001000101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101000001000010000100100001000101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100000010000100001001000010001010010100101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100000010000100001001000010001010010100101001010010100101001010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000000100001000010000100100010100101001010010100101001010010100101001010010000100011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000000100001000010000100100010100101001010010100101001010010100101001010010000100011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100110101101011010110101101011010001000010011100111001110011100111001110011100111001110011100010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001110011100100111001110011100111101011010111001110001010010100101001010010100101001010010100101001010111001110010011100111110011100111001110011100111001111111111111111111111111"),
                ("11111111111111111111111001110011100100111001110011100111101011010111001110001010010100101001010010100101001010010100101001010111001110010011100111110011100111001110011100111001111111111111111111111111"),
                ("11111111111110011100100111110011100100111001110011100111001110011111001110011100010100101001010010100101001010010100101000100111001110010011100111110011100100111001110011100111110011111111111111111111"),
                ("11111111111110011100100111110011100100111001110011100111001110011111001110011100010100101001010010100101001010010100101000100111001110010011100111110011100100111001110011100111110011111111111111111111"),
                ("11111111111110011100100111001110011111001110011100111001110011100111001110011111111001110011100111000010000100001000010000100001000010011100111001001110011110101101010011100111001111100111001111111111"),
                ("11111111111110011100100111001110011111001110011100111001110011100111001110011111111001110011100111000010000100001000010000100001000010011100111001001110011110101101010011100111001111100111001111111111"),
                ("11111111111110011100100111001110011100111001110011100111110011100111111111111111111111111111111111111110011100001000010000100001000010000100001001001110011100111001110011100111101011100111001111111111"),
                ("11111111111110011100100111001110011100111001110011100111110011100111111111111111111111111111111111111110011100001000010000100001000010000100001001001110011100111001110011100111101011100111001111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011111111111111111111111111111111111111001110000100001000010000100001001001110011100111001110011100111101011100111001111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011111111111111111111111111111111111111111111111100001000010010011100111001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111001110011111001110011111111111111111111111111111111111111111111111100001000010010011100111001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111001110010011100111001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001001110011110101101011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001001110011110101101011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_R_4.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111101011010110101101010011100111110011100111111111111100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111101011010110101101010011100111110011100111111111111100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111001110011100111001110011100111110011100111001110000100000010000100001000010010000100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001100001000010010000100000010000100001000010000100001000010000100001000010000100100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001100001000010010000100000010000100001000010000100001000010000100001000010000100100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111101111011110111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111000010000110111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111000010000110111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000110111101111011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000110111101111011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010100101001000010000001000010000100001000010100101001010010100101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010100101001000010000001000010000100001000010100101001010010100101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000101001000010000100001000010100101010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000101001000010000100001000010100101010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000100000010000100001000010101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000100000010000100001000010101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101001010001000010000001000010000100001010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011100111001110011100010100101001010010100101000100001000000100001000010000101000111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011100111001110011100010100101001010010100101000100001000000100001000010000101000111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001111100111000010000100111001110011100111001110011100111000010000100110101101011010110101101011100111001111111111111111111111100111001110011111111111111111111"),
                ("11111111111111111111111001001110011100111001111100111000010000100111001110011100111001110011100111000010000100110101101011010110101101011100111001111111111111111111111100111001110011111111111111111111"),
                ("11111111111111111111111001001110011111001110000100001000010000100001000010001010010100101001010010100101001010100111001110011110101101011100111001111111111111001110010011100111001111100111001111111111"),
                ("11111111111111111111111001001110011111001110000100001000010000100001000010001010010100101001010010100101001010100111001110011110101101011100111001111111111111001110010011100111001111100111001111111111"),
                ("11111111111110011100111001110011100001000010000100001000010000100001000010001010010100101001010010100101001010100111001110011100111001111100111001110011100111001110010011100111001110011100111110011100"),
                ("11111111111110011100111001110011100001000010000100001000010000100001000010001010010100101001010010100101001010100111001110011100111001111100111001110011100111001110010011100111001110011100111110011100"),
                ("11100111001101011010100110010000100001000010000100001000010000100111001110011100111001110011100111001110011100111001110011100111001110000101001010010100101100111001110011100111001110011100111110011100"),
                ("11100111001101011010100111001110011001000010000100001001110011100111111111111111111111111111111111111111111111111111111111100001010010100101001010010100101100111001110011100111001110011100111110011100"),
                ("11100111001101011010100111001110011001000010000100001001110011100111111111111111111111111111111111111111111111111111111111100001010010100101001010010100101100111001110011100111001110011100111110011100"),
                ("11100111001101011010100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111001110000101001011001110011100111001110011100111001111100111001111111111"),
                ("11100111001101011010100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111001110000101001011001110011100111001110011100111001111100111001111111111"),
                ("11111111111110011100110101001110011100111001111010110101110011100111111111111111111111111111111111111111111111111111111111111111111111111100111001001110011100111001110011100111001111100111001111111111"),
                ("11111111111110011100110101001110011100111001111010110101110011100111111111111111111111111111111111111111111111111111111111111111111111111100111001001110011100111001110011100111001111100111001111111111"),
                ("11111111111110011100110101001110011100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100100111001110011100111110011111111111111111111"),
                ("11111111111110011100110101001110011100111001110011100111110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100100111001110011100111110011111111111111111111"),
                ("11111111111111111111111001101011010100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_R_5.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111101011010110101101010011100111110011100111111111111100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111101011010110101101010011100111110011100111111111111100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111001110011100111001110011100111110011100111001110000100000010000100001000010010000100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111110011100100111001110011100111001110011100111110011100111001110000100000010000100001000010010000100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111001001110011100111001100001000010010000100000010000100001000010000100001000010000100001000010000100100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000011011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111101111011110111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111101111011110111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111000010000110111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000000100001000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111000010000100000010000100001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000110111101111011110111101111011110111111001110010111101111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000110111101111011110111101111011110111101111011101001010011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010100101001000010000001000010000100001000010100101001010010100101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010100101001000010000001000010000100001000010100101001010010100101001010010100111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000101001000010000100001000010100101010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000101001000010000100001000010100101010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000100000010000101010010100101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000100000010000101010010100101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000100000010000101010010100101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000101001010010100101000100000010000101010010100101001010010100101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010001000010000001000010101001010010100101001000111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000101001010111001110011100001000010011010110101101011010110101101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011100111000101001010111001110011100001000010011010110101101011010110101101001010111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100010100101001010010100101010011100111001110011110101101011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100010100101001010010100101010011100111001110011110101101011100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100001000010001010010100101010011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100001000010001010010100101010011100111001110011100111001111100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100001000010000100111001110011100111001110011100111001110000101111001110011111111111110011100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100001000010000100111001110011100111001110011100111001110000101111001110011111111111110011100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000010000100001000010000100111001110011100111000010100101001010010100101001010010111100111001001110011100111001111100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011001000010000100111001110011111111111110011100001010010100101001010010110011100111001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011001000010000100111001110011111111111110011100001010010100101001010010110011100111001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111001110011100111001110011111001110011100111001111111111111001110000101100111001110011100111001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111111110011100100111001110011100111001110011100111001110011111001110011100111001111111111111001110000101100111001110011100111001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111111110011100110101101010011100111001110011100111001110011110101101010011100111110011100111001110010011100111001110011100111001110011100111001111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100110101101010011100111001110011100111001110011110101101010011100111110011100111001110010011100111001110011100111001110011100111001111100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101101011010100111001110011100111001110011100111110011100111001110010011100111001110011100111110011100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101101011010100111001110011100111001110011100111110011100111001110010011100111001110011100111110011100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100110101101011010100111001111100111001111111111111111111111100111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_U_0.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000001000010010000100010100101011100111001110011100111001110011100111001110011100010100101000100001000000100001111001110011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100111001110000001000010010000100010100101011100111001110011100111001110011100111001110011100010100101000100001000000100001111001110011100111001111111111111111111111111"),
                ("11111111111111111111111001101011010110101101011010110101110011100010100101001010010100101001010010100101001010010100101001010010100101011100111001101011010110101101011010110101110011111111111111111111"),
                ("11111111111111111111111001101011010110101101011010110101110011100010100101001010010100101001010010100101001010010100101001010010100101011100111001101011010110101101011010110101110011111111111111111111"),
                ("11111111111111111111111001101011010100111001110011100111110011100001000010001010010100101001010010100101001010010100101001010001000010011100111001001110011100111001111010110101110011111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111110011100001000010000100111001110011100111001110011100111001110000100001000010011100111001001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111001001110011100111001110011100111110011100001000010000100111001110011100111001110011100111001110000100001000010011100111001001110011100111001110011100111110011111111111111111111"),
                ("11111111111111111111111111110011100111001110011100111001110011100001000010000100111001110011111111111111111111111001110000100001000010011100111001110011100111001110011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100111001110011100111001110011100001000010000100111001110011111111111111111111111001110000100001000010011100111001110011100111001110011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011111111111111111111111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011111111111111111111111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010100111001110011111001110011111111111111111111111001110010011100111001111010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010100111001110011111001110011111111111111111111111001110010011100111001111010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011111001110011111111111111111111111001110010011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011100111001111010111001110011111111111111111111111001110011010100111001110011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011100111001111010111001110011111111111111111111111001110011010100111001110011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010110101101011100111111111111111111111111111111111111111111100110101101011010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010110101101011100111111111111111111111111111111111111111111100110101101011010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110011111111111111111111111111111111111111111111111111111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_U_1.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010001010010100100001000010000100001010010101010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000000100001010100101001010010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100010100101001010010100101001010010100101001010010100101001010010100101011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100010100101001010010100101001010010100101001010010100101001010010100101011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010010000100111001110001010010100101001010010100101001010010100101001010111001110011100111000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101101011010110101101011100111001110011100111001110011100111001110011100010100101011100111001101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101101011010110101101011100111001110011100111001110011100111001110011100010100101011100111001101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011110101101001010010100101001010010100101001010010100101001010111001110010011100111101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001100100010100101001010010100101001010001000010000100111001110010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001100100010100101001010010100101001010001000010000100111001110010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100001000010000100111001110011100111001110011100001000010000100111001110011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100001000010000100111001110011100111001110011100001000010000100111001110011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100001000010011100111000010000100100111001111010100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100001000010011100111000010000100100111001111010100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001100100001000010011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001100100001000010011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010100111001110011110101101011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011110101101011010110101101010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011110101101011010110101101010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_U_2.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010110101101011010100111001101010010100101001010010100101001010010100101011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111101011010110101101011010100111001101010010100101001010010100101001010010100101011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011110101101010011100111001101010010100101001010010100101001010111001110011100111001001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001111100111001110011100111001110011100010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011100111001110011100111001111100111001110011100111001110011100010100101011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011010100101001010010100101001010010100101001010111001110011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100001000010011100010100101001010010100101001010100111001111010100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100001000010011100010100101001010010100101001010100111001111010100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011001000010000100111001110011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001101011010100111001100100111001110011100111001001110011110101101011010110101101010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101011010111001110011100111001001110011100111001110011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111111111111111111111110011100100111001110011100111001111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_U_4.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100010100101001010001010010100100001000010000100001010010101010010100101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100010100101001010010100101001010010100101001010100111001111010110101101011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100010100101001010010100101001010010100101001010100111001111010110101101011010110101001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111110011100111001110001010010100101001010010100101001010100111001110011110101101010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101011100111001110011100111001110011100100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101011100111001110011100111001110011100100111001110011100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100111001110001010010100101001010010100101001010010100101010011100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101010011100111001101010010100101001010010100101011100001000010000100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100110101101010011100111001101010010100101001010010100101011100001000010000100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100111001110000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011110101101011010110101101010011100111110011100111001110000100100111001111010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- character_U_5.bmp
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100001000010000001000010000100001001000010011100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001000010000001000010000110011100111001110011000010000100001001000010011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001100111001111010110101101011010100111001100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001100111001110011100111001110011100111001100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000010000100001000010000100001000010000110011100111001110011000010000100001000010000100001000010000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111100111001111111111111111111111111"),
                ("11111111111111111111111111110011100001000010000001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010011100111001111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010000100111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111000010000100000010000100001000010000100001000010000100001000010000100001000010000100100001001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100001010010100100000010000100001000010000100001000010000100100001010010111100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010001010010100100001000010000100001010010101010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100010100101001010010100101001010010100101001010010100101001010010100101000001000011110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100010100101001010010100101001010010100101001010010100101001010010100101000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100010100101001010010100101001010010100101001010010100101001010010100101000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110000001000011110011100111001110001010010100101001010010100101001010010100101001010111001110000100001000000100001111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101110011100010100101011100111001110011100111001110011100111001110011100110101101011010110101101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101110011100010100101011100111001110011100111001110011100111001110011100110101101011010110101101011010111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110011010110101001110011111001110001010010100101001010010100101001010010100101001010110101101010011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011111001110000100001000010001010010100101001010010100101000100100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111001110010011100111001110011111001110000100001000010001010010100101001010010100101000100100111001110011100111001110011111001110011111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100111001110000100001000010011100111001110011100111001110000100001000010011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001110011100111001110000100001000010011100111001110011100111001110000100001000010011100111001110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001111010100111001100100001001110011100001000010000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001111010100111001100100001001110011100001000010000100001000010010011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100001000010000100100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100001000010000100100111001110011100111110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011100111001110011100111001110011100111110011100110101101010011100111001111010110101110011100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011110101101011010110101101010011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111100111001001110011110101101011010110101101010011100111110011100111001110011010110101101011100111001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111110011100100111001110011100111001111100111001111111111111111111111100111001110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_0-0.png
                ("11111111111111111111111110110011001110011100110110110100100101001010010100111000101101001110011010010100101001100111001110011101101001111001110011100111001110011100111001111011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001100111101011000110001100011000100111011010110110100100101001110101101011010100111011011001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011011010011100111001110110101101001110011010010100111000110001100011000100111011010011100111001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011011010011100111001110110101101001110011010010100111000110001100011000100111011010011100111001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111011001100111001110011100111001100111011010110101101011010011110100100101001010010100101001010010100111010101101011010110101101100111001110011100111001110011100111111111111111111111"),
                ("11110111101111011110011001100111001110011100110011101101011010110101101011011010010011101011010110100100111010110101101011010100111001111001110011100111001110011100111001110011100101100011000110011001"),
                ("01110011100110001100110011100111001110011100110011101101011010110101101011011010010011100011000010010100111000110101101010011101101100111001110011011010011100111100111001110011100111001100111001101100"),
                ("01110011100110001100110011100111001110011100110011101101011010110101101011011010010011100011000010010100111000110101101010011101101100111001110011011010011100111100111001110011100111001100111001101100"),
                ("11101011001100111001100111100111001110011100110011110011001111001110011001111000110101101011010010010100101001100111001110110101101001111001110011011010110110011100111001110011100110011100111001101100"),
                ("11001110011100111001100111011011001110011001110011110011100111001110011001111000110101001110011110100100101001110101101011010100111001110011100111100110011100111100111001110011001110110110011100111001"),
                ("11001110011100111001110011100110011100111011010110101101001111001110011001111000110001101011010110000100101001110001100001001110101011010110101101001110011101101001110011100111100111001110011100110011"),
                ("11001110011100111001110011011010110101101011010110100111001110011100111101001001010010100101001010010100101001010010100101001110101011010011100111011010110101101011010110101101001110011100111001110110"),
                ("11010110101001110011100111011010110101101011010110110101100010011100111101011010110000100101001010010100101001010010100101001010011100010011100111011010110101101011010110101101011010110101101011010110"),
                ("11010110101001110011100111011010110101101011010110110101100010011100111101011010110000100101001010010100101001010010100101001010011100010011100111011010110101101011010110101101011010110101101011010110"),
                ("01001110001001110011101101011010110101101011010011110101011010011100110100101001110101101011010010011100001001010010100101001010011101010011100111011010110101101011010110100111001110011101101011010110"),
                ("01001110101001110011101101001110110101101011010011110101011010110101101101001001110000100001000010010100101001010010100101001110001001110011100111011010011101101001110011110001100011000110101101001100"),
                ("01001110101001110011100111001110011100111011010110110001101010110101101001111000010010100001000010000100101001010010100101001110001001111010110101101011010101101001110011110000100101001010010100111110"),
                ("01001110101011010110101101011010011100111001110011110001100011010110101101011010010010100001000010010100101001010010100101001110000100101000010000100111000010011101011010110100100101001010010100111010"),
                ("01001110101011010110101101011010011100111001110011110001100011010110101101011010010010100001000010010100101001010010100101001110000100101000010000100111000010011101011010110100100101001010010100111010"),
                ("01001010011001110011101101011010011100110100101001110001100001001010010100111000010010100101001110000100101000010010100111000010010100001000010000100101001010011101011010110100100111000010010100111000"),
                ("11000110000100101001010000100010011100111100001001010010100101001010010100101001110001100011000010010100101000010010100101001110001101001001010010100101001110101101011010010011101011000010010100101001"),
                ("01001010010100101001010000100101000010000100111000010010100001001010011101001001110000100101001010000100001001010010100101001100111001111010110101101010011100111101011010110001001111010110101101001001"),
                ("01001010010100101001110001101001001010011101011000010010100110011100111001101001110000100101001010000100001000010010100101000010011101010011100111001110011101101001110011100111001101001110001100001001"),
                ("01001010010100101001110001101001001010011101011000010010100110011100111001101001110000100101001010000100001000010010100101000010011101010011100111001110011101101001110011100111001101001110001100001001"),
                ("11000010011101011010100111011010110101101001101001010010100111010110101001101001010010100101001010010100001001010010100101001010010100111000110001001111000100111011010110101101001110011010010100111010"),
                ("01001010011101011010101101011010110101101001110011100111101011010110101101011000010010100101001010010100111000010010100111000010010100101001010011101010011101101011010110101101100111001100111001111000"),
                ("11010100111011010110101101011010110101101011010110101101011010110101101001101001010010100101001010010100101001010010100101001010011101011010110101001110110101101011010110100111100110110100111001111010"),
                ("10011101101011010110110011001110110101101011010110101101011010110101101011011010110101100011000010010100101001010010100111010100111011010110101101011010110101101001110011110011001110011100111001110011"),
                ("10011101101011010110110011001110110101101011010110101101011010110101101011011010110101100011000010010100101001010010100111010100111011010110101101011010110101101001110011110011001110011100111001110011"),
                ("11001110011011010110100111100110011100111011010011101101011010011100111011010110100110100101001110001101011010010010100110011101101011010110101101001110110100111100111001110011011010011100111001110110"),
                ("01100110011100111001110011100111001110011100111001110011100111001110011100110011110000100101001110001011010110100111001110011110011001110110101101011010011110011100111001110011100110011100111001111110"),
                ("01110111011100111001110011100111001110011100111001110011100111001110011100110011010011100011000110101001110011100111001111010110011100110011100111100111001110011100111001110011100111001110011100101100"),
                ("11110111011100111001110011100111001110011100111001100111001111001110011100111010010010100101001110001101011010110101101011000100111011010110101101100111001110011100111001110011100111001110011100111001"),
                ("11110111011100111001110011100111001110011100111001100111001111001110011100111010010010100101001110001101011010110101101011000100111011010110101101100111001110011100111001110011100111001110011100111001"),
                ("11001110011100111001011001100111001110011100111001110011011010110101101011010110110100100101001010010100101001010010100111010101101011010011100111100111001110011100111001110011100111001011000110001100"),
                ("11111111111111111111011001100111001110011100111001110011011010110101101011010110100110100101001010010100101001110101101010011101101011010110101101100111001110011100111001110011100111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011011010110101101011010110100111001110011110000100001000100111001110011100111001111001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111011001110011100111001110011011010110101101011010110101101011010110100111100001001110101101010011100111100111001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111011001110011100111001110011011010110101101011010110101101011010110100111100001001110101101010011100111100111001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111100110001100011001100111001100111100110011100111101010011100111011010110110100100001001010000100001000010011001111001110011100111001110011100111001110011001111111111111111111111"),

                -- explosion_0-1.png
                ("11111111111111111111111111111111111111111111001100110011011010011100110100101001110000100101001010010100101000110101101010011101101100110110101101001111001110011100111001111101111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011011010011100111100001001010010100101001010010100101001110001100010011101101100110011100111001111001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111110110011001110011100110011101101011010110101101001111010100111101011010110000100101001110101101010110101101001110110101101001111001110010110001100111111111111111111111111111111"),
                ("11111111111111111111111110110011001110011100110011101101011010110101101001111010100111101011010110000100101001110101101010110101101001110110101101001111001110010110001100111111111111111111111111111111"),
                ("11111111111111111111111110110011001110011100110011101101001110011100111011010110101101011010110110001101011000100111001110011101101001111001110011001110110110010110001100111111111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001101101001111010110101101011010110101011010110010010100110011100111001110011101101100111001110011100111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111110111001100011001001110110101101011010011100111001110011110001101011010010000100110011100111001110110101101001111001110011100111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111110111001100011001001110110101101011010011100111001110011110001101011010010000100110011100111001110110101101001111001110011100111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111110111001100011001001110110100111011010110101101011010110110100100001000010000100001001100111001110110101101100111001110011100111001110011100111001111101111111111111111111111111"),
                ("11111111111111111111111110111001100011001011011001110011011010110101101011010011010010100001000010000100111010101101011010011100111100110011100111001111001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111111111101100011001100111001100111011010110101101011011010010010100101001010011100010011101101011010011100111100110110101101001111001111101111011110111111111111111111111111111111"),
                ("11111111111111111111111111111111001110011001110110101101011010110101101001110011100110100101001010010100110011101101011010011101101011010011100111100111001011001111011110111111111111111111111111111111"),
                ("11111111111111111111111111011011001110011100111001101101011010011100110100111000110101100011000010010100011010100111001110011101101011010011100110110011001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111111011011001110011100111001101101011010011100110100111000110101100011000010010100011010100111001110011101101011010011100110110011001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001100111011011010110100100101001110101101011010110100100101001110001100010011110011001110011100111100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111100111001110011011010110100111001110011100110100111000010011100011000110100100101001010010100111010101101100111001110011011010110101101001110011100111111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001101101011010011100111001110011100111101011010010010100101001110001100010011101101001111001110011011010110101101100111001110011111111111111111111111111"),
                ("11111111111111111111111111111011001110011100111001100111011010110101101001110011110101100011000010010100101001010010100110011101101011011001110011001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111011001110011100111001100111011010110101101001110011110101100011000010010100101001010010100110011101101011011001110011001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011011010110101101011010110110000100101001010010100101001010010100101001101101001111001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011001110011100111001111010110000100101001110001100011000010010100101000100111011011001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011100111001110011100101001010010100101001010010100111000010000100001001100111100111001110011100111001011001100111001011001111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011100111001110011011010011110101100011000010010100101001010010100101001110101001111001110011100111001011000110001100111111111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011100111001110011011010011110101100011000010010100101001010010100101001110101001111001110011100111001011000110001100111111111111111111111111111111"),
                ("11111111111111111111111111111001100011001100111001100111011010011100111101010011101101100011000010010100101001110001100001001110101011010011100111100111001011000110001100111111111111111111111111111111"),
                ("11111111111111111111111111111001100011001100111001101101011010011100111101010011101101100011000010011100011000010010100110011101101001110011100111001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111011001110011100110011101101011010011100111101010011101101100011000110101001111010110101101010110101101011011001110011001111001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111110110011001110011100110011101101011010110101101001110011100110100101001110101001111010101101011010110101101011010011100111100111001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111110110011001110011100110011101101011010110101101001110011100110100101001110101001111010101101011010110101101011010011100111100111001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111110110011101111010110011001100111011010110101101001110110110100100001000010011101010011100111001110110101101011011001110011100111001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111111111101100011001001111001110011001110110101101011010011110000100101001010010100101001110001100010011101101011011001110011100111001011001111011110111111111111111111111111111111"),
                ("11111111111111111111111111111111001110011001111001110011100110110101101011010011110101101011010110000100101000010010100110110101101011011001110011100111001111100110001100111111111111111111111111111111"),
                ("11111111111111111111111111110111001110011001110011110011100110110101101011010110101101101011010010010100101000010000100010011100111011011001110011100111001011001100111001110011111111111111111111111111"),
                ("11111111111111111111111111110111001110011001110011110011100110110101101011010110101101101011010010010100101000010000100010011100111011011001110011100111001011001100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100110011100111001110110101101011010011110100100101001110100100101001010010100111010101101011010011100111100110011110010110001100111101111111111111111111111111"),
                ("11111111111111111111111111100111001110011100110011101101011010110101101011010011010011101011010100111101001001110001100010011101101011011001110011100110110100111100111001111101111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001101101011010110101101011010110110101101011010100111001101001110001100010011100111001111001110011100110110101101100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001100111011010011100111001110110100111001110011100111100011000100111001110110101101011011001110011100110110101101100111001110011111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001100111011010011100111001110110100111001110011100111100011000100111001110110101101011011001110011100110110101101100111001110011111111111111111111111111"),
                ("11111111111111111111011001100111001110011100111001101101011011010110100100110011100111101011010110101001110011100111001110011100111001111001110011100111001100111100111001110011100111111111111111111111"),

                -- explosion_0-2.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("01100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11001110011100111001110010110011101111011111111111011000110011110111101111011110011001111111111111110110011110110011100111001110011011011111111111111101110011100111001110011000110001100111111111111111"),
                ("11001110011100111001110011100111001110011100101100111011100111001110010110001100110011100111001110011100111001110011100111001110011100111001110010110001100011000110001100110011100111001110011100111111"),
                ("11001110011100111001110011100111001110011100101100111011100111001110010110001100110011100111001110011100111001110011100111001110011100111001110010110001100011000110001100110011100111001110011100111111"),
                ("11001110011100111001110011100110011100111001110011011001100111001110011100111001110011100111001110011100111001110011100110110110011100110011100111100110110100111001110011110011100111001110011100111110"),
                ("11001110011100111001100111001110011100111100111001110011001110011100111100111001110011100111001110011100111001110011100110110110011100110110101101100111001101101011010110110011001110011110011100101100"),
                ("10110100111011010110101101001111001110011100111001100111011010110101101011010011110011100111001110011100110011101101011010011100111011010110101101001111001100111011010110101101011010110110011100111001"),
                ("10110101101011010110101101001111001110011100110011101101011010110101101011010110110011100111001100111011010110101101011010011101101011010110101101011010110101101011010110100111001110110101101011010110"),
                ("11010100111011010110101101011010110101101011010110101101011010011100111001110011110011100111001100111011010110100111001110011110101001110110101101011010110101101001110011110101001110110100111001110011"),
                ("11010100111011010110101101011010110101101011010110101101011010011100111001110011110011100111001100111011010110100111001110011110101001110110101101011010110101101001110011110101001110110100111001110011"),
                ("01001100111011010110101101011010110101101011010110100111001111010110101101011010101101100111001100111011010011100111001101001010010100110011100111011010110101101001110011110101011010011110001100001001"),
                ("10011101101011010110100111001110110101101001110011101101001110011100111001110011100110100101001110101011010011100111001111000010011100010011100111101010011101101001110011110101011011010010010100101001"),
                ("10011100111101011010010011101010110101101101011000110101001110110101101011010110110100100101001110001100011010100111001101001110101101010011100110100101001110101100011000110101011010011010010100111000"),
                ("11010100111101011010110100100111010110101101001001010000100111000110001100011000110000100101001010010100111000110101101011000110101100001001010010100101000010001101011010101101011011010010010100101001"),
                ("11010100111101011010110100100111010110101101001001010000100111000110001100011000110000100101001010010100111000110101101011000110101100001001010010100101000010001101011010101101011011010010010100101001"),
                ("11010100111001110011100111101001001010011100001001010011101011010110100100101001010010100101001110000100101001010010100111010110100100101001010010100101000010000100001000010011100011000010010100101001"),
                ("10011110001001110011110100100101001010010100101001110101001110011100111100001001010010100101001110000100101001010010100101001010010100001001010011100001001010000100101001010011101001001010010100101001"),
                ("10011110000100101001010010100101000010000100001001100111101011010110101100001001010011100011000110000100101001010010100101001010011101010011100111001111010010011001110011100111100001001010010100101000"),
                ("10011100111100011000110000100101000010000100111000100111011011010110100100111000010010100001000010010100101001110001100001001110001001110110101101011010110100111001110011100111001111010110001100011010"),
                ("10011100111100011000110000100101000010000100111000100111011011010110100100111000010010100001000010010100101001110001100001001110001001110110101101011010110100111001110011100111001111010110001100011010"),
                ("10011101101001110011100111101010011100111011010011101101011010110101101001101001010010100101001010000100110011100111001111010100111001110011100111001110011101101011010110100111001110110100111001110011"),
                ("10011101101001110011101101011010011100111011010110101101011010110101101011011010110101001110011100111011010110101101011010110110011011010110101101001110011101101011010110101101011010110101101011010110"),
                ("10011101101001110011101101011010110101101011010110101101011010110101101001110110100111100111001101101001110110100111001111001100111011010110101101100111001110011001110011110011001110011110011100111001"),
                ("11001110011100111001110011001111001110011100111001110011001111001110011001110011110011100111001110011100111001110011100111001100111001110011100111011010011110011100111001110011100110110100111001110110"),
                ("11001110011100111001110011001111001110011100111001110011001111001110011001110011110011100111001110011100111001110011100111001100111001110011100111011010011110011100111001110011100110110100111001110110"),
                ("11001110011100111001110011100111001110011100111001110011100110011100111001111001110011100111001110011100110011101101011010110110010110011001110011001110011110011100111001110011001110011100111001110011"),
                ("11001101101011010110101101001111001110011100111001110011100111001110011100111001110011100111001110011100111001101101011010110110011100111001110011100111001110011100111001110011011011001110011100111001"),
                ("10011101101011010110100111100101100011001111001100110011100111001110011100101100011000110001100110011100111001101101011010110110011100101100011001111011001110011100111001110011100111001110011100111001"),
                ("11001110011100111001110010110011001110010110011110011000110011001110011100101100011001100111001110011100111001110011100110011110010110011110111101111001100110010110001100011000110001100011000110011001"),
                ("11001110011100111001110010110011001110010110011110011000110011001110011100101100011001100111001110011100111001110011100110011110010110011110111101111001100110010110001100011000110001100011000110011001"),
                ("11001110010110001100111101111011001110011111111111011101111001100011001100111111111110110001100110011100111001110011100110011110011111011111111111111101110111100110001100011001111111111111101111011110"),
                ("11001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_0-3.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111110011001100111001011001100111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111110011001100111001011001100111001110011100111001111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110010110011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111001110011100110011100111100111001110011100111001110011100111001100111001110011110011100111001110010110001100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111001110011100110011100111100111001110011100111001110011100111001100111001110011110011100111001110010110001100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011001110011100110110101101100111001110011100111001110011100111001100111001110011101101001111001110011100111001110011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111110110011001110011001111001110011100111001110011100111001110011100110110101101011010110101101001111001110011100111001110011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111100111001100111001111001110011001111001110011001110011110011100110110100111001110011100111100111001110011100111001110011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111101100011001100111001110011100110110101101100111001110011001110011100111001111001100111001111001100111001111001110011100111001110010110001100111111111111111111111111111111"),
                ("11111111111111111111111110110001100011001100111001110011100110011100111001111001110011011010110101101011010110101101011011001100111001110110101101011011001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111110110001100011001100111001110011100110011100111001111001110011011010110101101011010110101101011011001100111001110110101101011011001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011100110011100111001110110110011011010110101101011010110101101011010110101101011010110101101001111001110011100111001111011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011100111001110011001110110100111101011010100111011010011100111001110110101101011010110101101001111001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001100111100110011100111101010110110100100101001010011100001001100111001110110101101011010011100111100111001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011001110110101101001110110110100100101001110000100101001110101101010011101101001111001110011100111001110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011001110110101101001110110110100100101001110000100101001110101101010011101101001111001110011100111001110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011100110011100111011010011110000100101001010010100111010010010100101001110101001111001110011100111001110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011100111001110011011010011110000100101001010010100111010100111001111010110101001110011100111001111001110011100111001111011111111111111111111111111"),
                ("11111111111111111111111111111111001110011100110110100111100110110101101011010011010010100101001110101001110110101101011010110101101001110011100111011010110101101100111001111011111111111111111111111111"),
                ("11111111111111111111111111100111001110011001110110101101100110110101101011011010010010100101001110101001111010100111001110110100111101010011100111011010011100111100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011001110110101101100110110101101011011010010010100101001110101001111010100111001110110100111101010011100111011010011100111100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011001110110101101011010110101101011010011110100100101001100111101011000110101101010011100111011010011100111100111001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011100110110101101011010110101101011011010110101101011010100111101010011110101101001001100111011011001110011100111001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001101101011010110101101011010011110001001110011100111101010011100111001110011101101011010011100111100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111111110111101100111001110011011010110101101011010110100111001110011110000100101001100111001110011100111011010110101101100111001110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111111111110111101100111001110011011010110101101011010110100111001110011110000100101001100111001110011100111011010110101101100111001110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111111101110011101111001100110011100110011100111011010110101101100011000010010100111000100111001110011100111011010110101101100111001110010110001100111111111111111111111111111111"),
                ("11111111111111111111111111111011110111101111011110110011100110011100111011010110100110100101001010010100111000100111001111010100111001110011100111011010011110011110111101111101111111111111111111111111"),
                ("11111111111111111111111111111011110111101100111001110011001110011100111011010011110000100101001010011101011010110101101010011100111001110011100111011010110110011111011110111101111111111111111111111111"),
                ("11111111111111111111111111111001100011001100111001100111011010011100111011010110110100100101001110001101011000110001100011010100111001110011100111001111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111111111001100011001100111001100111011010011100111011010110110100100101001110001101011000110001100011010100111001110011100111001111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111110111001100011001100111001100111011010110101101001110011100111101011010110001101011010110101101011010110101101010011100111001110011110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110111001100011000110011001100111011010011100111101010011101101101011010010011101011010110001100011000110101101010011100111001110011011001111011110111011111111111111111111111111"),
                ("11111111111111111111111101111011110111101100111001110011011010110101101001110110100111100011000010010100111010100111001111010110101100011010110101001110011110010110001100011001111111111111111111111111"),
                ("11111111111111111111111110111001100011001100111001100111001110011100111001110110100111101011010010011100011010110101101011010100111101011010110101001110011110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110111001100011001100111001100111001110011100111001110110100111101011010010011100011010110101101011010100111101011010110101001110011110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110111001100011001100111001110010110010011100111001110011100111101011010110101100011010110101101010011100111001110011100111001111001111101111011110111011111111111111111111111111"),

                -- explosion_0-4.png
                ("11111111111111111111111111110111110111101111011001100111001110011100111001110011110101101011010110001101011010100111001110011100111001101100011001100111001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111111100111001110011100110011100111101011010110101001111010110101101011010110000100111010100111001110110100111001110011100111001111001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111110110001100011001100110011100111101011000110001101011010100111101011010010010100111000100111001110110100111011010110101101100111001110011111011110111101111011111111111111111111"),
                ("11111111111111111111111110110001100011001100110011100111101011000110001101011010100111101011010010010100111000100111001110110100111011010110101101100111001110011111011110111101111011111111111111111111"),
                ("11111111111111111111111111110111110111100110010011100111001111010110101101011000110001101011010110100100111010101101011010011110101001110110101101001111001011000110001100011101111111111111111111111111"),
                ("11111111111111111111111111100111001110011100110011100111001111010110101101011010110101101011010110101100011010100111001110011100111011010110101101001111001110010110001100011101111111111111111111111111"),
                ("11111111111111111111111110110001100011001100111001100111001110011100111001111010110001100011000110101100001001110101101010110101101001110110101101001111001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111110110001100011001100111001100111001110011100111001111010110001100011000110101100001001110101101010110101101001110110101101001111001110010110001100111101111111111111111111111111"),
                ("11111111111111111111111111111011110111101100110110101101001110011100111001110011110101101011010110100100101001110001100010011101101001110011100111100111001110011111011110111101111111111111111111111111"),
                ("11111111111111111111111111111011101111011100110011101101001110011100111001111010100111100011000010010100101001100111001110110101101001111001110011100111110111101111011110111101111111111111111111111111"),
                ("11111111111111111111111111111101100011001100111001110011011010110101101001110011100111100011000010010100111000101101011010110101101001111001110011100101100111100111001110111111111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011011010110101101001110011100110100101001010011100010011100111001110110101101011010110101101100111001110011111011110111111111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011001110110101101011010011100111001110011110101001110011110001100010011101101011010110101101011011001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011100111001110011001110110101101011010011100111001110011110101001110011110001100010011101101011010110101101011011001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011100110110101101001101001110101001110011110101001111010110101101011010101101011010110101101011010110110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011001110110101101001110011110101100011000110101001101001110101101010011101101011010110101101011010110100111100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011001110011101101001111010110101001110110100111101011010100111101001001010010100111010101101011011001110011011010110100111100111001110011111111111111111111111111"),
                ("11111111111111111111111111110111001110011011010110101101001110011100111011010110101101011010110100111101001001010010100110011101101011011001110011001110110110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111110111001110011011010110101101001110011100111011010110101101011010110100111101001001010010100110011101101011011001110011001110110110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111110111001110011100111001100111001110011100111101011010100111101011010010010100101001110001100010011101101100111001110011100111001110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011100110011100111101001001010011101011010010010100101001110001100010011101101001111001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111111111111001110011100111001110011100110011100111011010011110100100101001010011100001001110101101010110100111011010011100111100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011001110110101101011010110100110100101001110000100101001110101101010110110101001111001110011001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001110011001110110101101011010110100110100101001110000100101001110101101010110110101001111001110011001111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110110011001110011100111001100111011010110101101011010110100111001110011101101001111010100111001110110100111100111001110011100111001110011100111001011001111111111111111111111111"),
                ("11111111111111111111111111110111001110011100111001100111011010110101101011010110101101011010110101101011010110110011100110110100111001111001110011100111001110011100111001110011111111111111111111111111"),
                ("11111111111111111111111110111001100011001100111001101101011010011100111001111001101101011010110101101011010110110011100111001100111001111001110011100111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111111111101100011001100111001110011100110011100111001111001100111100111001100111001110011110011100111001110011011011001110011100111001110010110001100111111111111111111111111111111"),
                ("11111111111111111111111111111101100011001100111001110011100110011100111001111001100111100111001100111001110011110011100111001110011011011001110011100111001110010110001100111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111100111001110011100111001110011001110011100111011010110110011100110011110011100111001100111100110011100111001111001110011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111100111001110011100110011100111011010110101101011010110110011100111001110011100111001110011100110011100111100111001011001111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111100111001110011100110011100111011010011100111100111001110011100111001110011100111001110011011011001110011100111001111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111101100011001100111001110011100110011100111100111001110011100111001110011100111001110011001111001110011100111001111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111101100011001100111001110011100110011100111100111001110011100111001110011100111001110011001111001110011100111001111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111011001100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110010110011001011000110011110111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_0-5.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("01110011101111011110011100111011110111101111011110111111111101100011001100111001110011111111111111111100111001110011100101100110010110011111111111111111111111111111111111111111111111111111111111111111"),
                ("01100011001111011110011000110001100011001111011110011101111011001110011100111001110011100111001110011100111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111"),
                ("01100011001111011110011000110001100011001111011110011101111011001110011100111001110011100111001110011100111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111"),
                ("11001110011100111001011001100111001110011100111110111101100111001110011100110011100111100111001110011100111001110011100111001110011100111001110011100101100111101111111111111111111111111111111111111111"),
                ("11001110011100111001110011100111001110011100111110011001100111001110011011010110101101011010110110011100111001110011100111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("11001100111100111001100111001110011100111100111001110011100110110101101011010110101101001110011110011100111001100111001111001110011100111001110011001111001110011100111001110011111111111111111111111111"),
                ("01100100111011010110101101011010110101101001111001110011011010110101101011010110110011100111001110011100110011110011100111001110011100111001110011001110011110011100111001110011111111111111111111111111"),
                ("10011100111011010110100111011010011100111001110011100111011010110101101011010110101101011010110110011001110110100111001111001100111001110110101101100111001101101001110011110011111111111111111111111111"),
                ("10011100111011010110100111011010011100111001110011100111011010110101101011010110101101011010110110011001110110100111001111001100111001110110101101100111001101101001110011110011111111111111111111111111"),
                ("10011100111001110011110101001110110101101011010110101101011010110101101011010110101101011010110101101011010011110101101010011100111001111001110011001111001110011100111001110011100111111111111111111111"),
                ("10011101101011010110100111001110110101101001110110101101011010011100111101010011110101001110011100111001110110101101011010110101101100111001110011100111001110011100111001110011100111110111111111111111"),
                ("10011100111001110011101101001111010110101100010011101101001111000110001101011010010010100101001110001100011010110101101010011110011100111001110011100111001110011100111001110011100101100111111111111111"),
                ("11010110101100011000110101101001001010010100101001110001001110011100111101001001010010100101001010010100101001010010100111010101101011010011100111001111001110011100111001110011100111001111111111111111"),
                ("11010110101100011000110101101001001010010100101001110001001110011100111101001001010010100101001010010100101001010010100111010101101011010011100111001111001110011100111001110011100111001111111111111111"),
                ("11010010010100101001010011100011000110000100101001010011100010011100111001110011110101101011010010010100111000010010100110011101101011010011100111100111001110011100111001110011100101100111111111111111"),
                ("11000110000100101001110101101011010110101101001001010010100111010110101101011010100111001110011010010100101001110001100010110101101011010011100111100111001110011100111001110011100111001111111111111111"),
                ("11010110101101011010110101101011000110001101011000110000100110011100111001111000110101011010110110101101001001010010100110011101101011011001110011011010110110011100111001110011100111001111111111111111"),
                ("11010110101001110011110001101011000110001101010011100111001110011100111101011010100111011010110100110100111010100111001110011101101011010011100111001110110100111001110011110011100111001111111111111111"),
                ("11010110101001110011110001101011000110001101010011100111001110011100111101011010100111011010110100110100111010100111001110011101101011010011100111001110110100111001110011110011100111001111111111111111"),
                ("10011110101101011010110001101011010110101001111010100111001110011100110100110011101101011010110110100100110011101101011010110101101100111001110011001110110100111001110011110011100111001111111111111111"),
                ("10011100111101011010110101101010011100111001110011100111001110110101101001110011100111011010110110101101010110101101011010110101101001110011100111001110110101101100111001110011100111111111111111111111"),
                ("10011110101100011000110101101010011100111001110011101101011010110101101011010110110101001110011100111001110011101101011010110101101001110011100111100110011100111100111001110011111111111111111111111111"),
                ("10011110101101011010100111001110011100111001110011101101011010011100111100110011100111001110011100111100111001100111001110110101101011011001110011100111001110011100111001110011111111111111111111111111"),
                ("10011110101101011010100111001110011100111001110011101101011010011100111100110011100111001110011100111100111001100111001110110101101011011001110011100111001110011100111001110011111111111111111111111111"),
                ("10011100111001110011100111001110011100111011010110110011100111001110011100111001101101011010110100111100111001110011100110011100111011011001110011100111001110010110001100011001111111111111111111111111"),
                ("11001100111001110011100111001111001110011011010011110011100111001110011100111001100111011010110110011100111001110011100111001110011100111001110011100111001110010110001100111111111111111111111111111111"),
                ("11110110011100111001011001100111001110011100111001110011100111001110011100111001100111011010110110011100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("11110110010110001100111101100101100011001111011101011001100111001110011100111001110011100111001110011100111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111"),
                ("11110110010110001100111101100101100011001111011101011001100111001110011100111001110011100111001110011100111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111"),
                ("11101110010110001100111011100101100011001111011110111111111111001110010110001100011001110111101111011111111111011000110001100111010111011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_0-6.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111101110011101110101100011001111111111111111110111101011000110001100011001100111111111111111111110111100110001100110011110101100110011100111101"),
                ("11111111111111111111111111111111111111111111111111111110110001100011001100111001110011100111001110011100111001110011100111001110011100111001110010110011101111100110001100110011111001100110011100111110"),
                ("11111111111111111111111111111111111111111111111111111110110001100011001100111001110011100111001110011100111001110011100111001110011100111001110010110011101111100110001100110011111001100110011100111110"),
                ("11111111111111111111111111111111111111111100111001110011100111001110011100111001110011100111001110011100110110100111001111001110011100111001110011100111001110011100111001110010110011001110011100111110"),
                ("11111111111111111111111111111101100011001100111001110011100111001110011100111001110011100111001110011100110110100111001111001110011100111001110011100110011101101100111001100111001110011100111001111001"),
                ("11111111111111111111111110110001100011001100111001110011100110110101101001110011110011100111001110011001110110101101011011001110011100111001110011100110110101101001110011100111001110011100111001110011"),
                ("11111111111111111111111111100111001110011100111001110011100110110101101011010110100111100111001110011001110011100111001110011110011001110110101101011010011100111001110011100111001111010110101101010011"),
                ("11111111111111111111111111100111001110011001110011110011001110011100111011010110101101001110011100111001110011110101101010110101101011010110101101011010011100111001110011110101101011000110101101010011"),
                ("11111111111111111111111111100111001110011001110011110011001110011100111011010110101101001110011100111001110011110101101010110101101011010110101101011010011100111001110011110101101011000110101101010011"),
                ("11111111111111111111110011100111001110011011010110100111001110011100111011010110101101011010110110101101010110100111001110011100111011010011100111001110011100111001110011110101101011010100111001110011"),
                ("11111111111100111001110011100110011100111001110110100111100111001110011011010110101101001110011010011101010110101101011010011010011001110011100111001111010100111101011010110101100011010110101101010011"),
                ("11111111111100111001110011100110011100111001110110100111001110110101101011010011100111101011010010011001110110100111001111010110101001110011100111001110011110101100011000110101100010011110101101011010"),
                ("11111111111100111001110011100111001110011100110110101101100110110101101011010011010010100101001110101101010110110101101011000100111001101001010011100011000110101100011000110101101011010110101101011010"),
                ("11111111111100111001110011100111001110011100110110101101100110110101101011010011010010100101001110101101010110110101101011000100111001101001010011100011000110101100011000110101101011010110101101011010"),
                ("11111111111100111001110011100111001110011100111001110011001110110101101011010110110000100101001010010100110011100111001111010110101101001001010010100101001110101101011010110101101001001110001100011000"),
                ("11111111110110001100110011100111001110011100111001110011001110110101101011010011010011100011000010010100111010110101101010011100111001111000110000100101001010011100011000110000100101001010010100111010"),
                ("11111111111100111001110011100111001110011100111001100111001110110101101011011010010010100101001010010100101001010010100101001110101001110011100111100001001010010100101001110101101011000110101101011010"),
                ("11111111110110001100110011100111001110011100111001110011100111001110011100110011110101101011010110001100001001010010100111010110101100010011100111011010011110001101011010100111011010011100111001110011"),
                ("11111111110110001100110011100111001110011100111001110011100111001110011100110011110101101011010110001100001001010010100111010110101100010011100111011010011110001101011010100111011010011100111001110011"),
                ("11111111111111011110110011100111001110011100111001110011100111001110011011010110101101011010110100111001110011110101101010011110101001110110101101011010110100111011010110100111001110110101101011010011"),
                ("11111111111111111111110011100111001110011100111001100111100110011100111001110011110101001110011101101011010110101101011010110101101011010110101101011010110101101011010110100111101010011100111001110011"),
                ("11111111111111111111111111100110011100111011011001110011011010011100111001111001100111011010110100111100110110101101011010110101101011010110101101001110011100111001110011101101001110110100111001110011"),
                ("11111111111111111111111111100111001110011100110011100111100111001110011100111001110011001110011110011100111001110011100110110101101011010110101101100111001100111011010110101101011010110100111001101100"),
                ("11111111111111111111111111100111001110011100110011100111100111001110011100111001110011001110011110011100111001110011100110110101101011010110101101100111001100111011010110101101011010110100111001101100"),
                ("11111111111111111111111111100111001110011100111001100111100111001110011100111001100111100111001110011100110011101101011010110101101011011001110011100111001110011001110011100111001111001100111001111001"),
                ("11111111111111111111111111111111001110011100111001110011100111001110011100111001110011100111001110011100110110101101011010110101101100111001110010110011110110011100111001110011100111001110011100111001"),
                ("11111111111111111111111111111111111111111111001100110011100111001110011100111001110011100111001110011100111001100111001110011110011100111001110011111011110110011100111001110010110011001110011100111001"),
                ("11111111111111111111111111111111111111111111111111111110110001100011001100111001110011100111001110011100111001110011100111001110011100111110111100111011110111100110001100011000110011110011000110001100"),
                ("11111111111111111111111111111111111111111111111111111110110001100011001100111001110011100111001110011100111001110011100111001110011100111110111100111011110111100110001100011000110011110011000110001100"),
                ("11111111111111111111111111111111111111111111111111111111111101100011001100101100110011100111001110011111111111110011100111001110010110011111111111111111110111101111011110011100111011110011100111001110"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_1-0.png
                ("11001110011110111101111101100111001110011100111010010010100111000110000100101001010010100101001010000100001000010000100001000010011101011010110101101001001100111011010110101101001111001111101111011110"),
                ("11001110010110001100111011100110110101101001101001010010100101001010011100001001010000100001000010000100001000010010100101000010010100111000110000100111010100111001110011101101001111001011000110011001"),
                ("10011101101011010110100111001110011100111101001001110001100011000110001100001001010000100001000010000100001000010000100001001010000100111000110001101010011100111001110011101101011011001110011100101100"),
                ("10011101101011010110100111001110011100111101001001110001100011000110001100001001010000100001000010000100001000010000100001001010000100111000110001101010011100111001110011101101011011001110011100101100"),
                ("10110101101011010110101101011010011100111101011000010010100101001010010100101001010000100001000010000100001000010000100001001010010100111010110101101011000100111001110011101101001111001110011100111001"),
                ("10110101101011010110101101001110011100111001111010010010100101001010010100101000010000100001000010000100001000010000100001001010011100011010110100100111000100111001110011101101011010011100111001110011"),
                ("10110101101011010110101101101011010110101101001001010010100111000110000100101001010010100001000010000100001000010000100001000010011100011010110100100111000100111001110011101101011010110101101011010011"),
                ("10110101101011010110101101101011010110101101001001010010100111000110000100101001010010100001000010000100001000010000100001000010011100011010110100100111000100111001110011101101011010110101101011010011"),
                ("10011101101011010110101101001101001010010100101001010010100101001010011100001001010000100001000010000100001000010010100101001010010100101001010010100101001010011001110011101101001110110100111001110011"),
                ("01001100111011010110100111011011010110100100101001010010100101001010011100001001010000100001000010000100001001110001100001001010010100101001010010100101001010011101011010110100100111010110101101010011"),
                ("01001110101011010110110101101011000110000100101001110001100011000110001100001001010000100001000010000100001001110001100001001010011100011000110001100001001010010100101001010010100101001110101101010011"),
                ("11000110001101011010110000100101001010010100111000010010100101001010010100101000010000100001000010000100001001010010100101001010010100101001010010100111000010010100001000010011100011000010010100111000"),
                ("01001010010100101001010010100101001010010100101001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000010010100001000010010100001001110001100001001"),
                ("01001010010100101001010010100101001010010100101001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000010010100001000010010100001001110001100001001"),
                ("01001010010100101001110001100001001010010100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100001000010000100001001110001100001000"),
                ("01001010000100001000010010100101001010010100101000010000100101001010010100001000010000100001000010000100001000010000100001000010000100001000010001100001000010000100001000010000100111010010010100100011"),
                ("01001010000100001000010000100001000010000100101001010000100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010000100001000010000100001000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("01000010000100101001010010100101000010000100001000010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("01000010000100101001010010100001000010000100001001010011100001001010010100001000010000100001000010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100001001"),
                ("01000110001100011000010010100001000010000100101001010011100001001010010100001000010000100001000010000100001000010000100001001010000100101001010010100101001010010100001000010000100001000010000100001000"),
                ("01000110001100011000010010100001000010000100101001010011100001001010010100001000010000100001000010000100001000010000100001001010000100101001010010100101001010010100001000010000100001000010000100001000"),
                ("01001010010100101001010010100101001010010100001000010010100101001010010100001000010000100001000010000100001000010000100001000010010100101001010010100111000110000100101001010011100001001010010100101001"),
                ("01001010010100101001010010100101001010010100101000010000100101001010010100001000010000100001000010000100001000010000100001000010000100101001010010100001000010011100011000010010100111000110001100011000"),
                ("01001010010100101001110000100101001010010100101000010001100001001010010100101000010000100001000010000100001000010000100001000010000100111000110000100101000010011100011000010010100101001010010100101001"),
                ("11010110000100101001010010100111000110001100001001010011100011000110001100001001010000100001000010000100001000010000100001000010000100101000010001100001001010010100101001010010100101001010010100101001"),
                ("11010110000100101001010010100111000110001100001001010011100011000110001100001001010000100001000010000100001000010000100001000010000100101000010001100001001010010100101001010010100101001010010100101001"),
                ("11010110100100101001010011100001001010010100111000110000100101001010010100101001010000100001000010000100001000010000100001000010000100101000010000100111000010010100101001010010100111000100111001101001"),
                ("01001010011100011000010011101011000110000100101001010010100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010010100101001100111001111000"),
                ("11010110101001110011010011100010011100111100001001010010100111000110001100001001010010100101001010000100001000010000100001000010010100101000010000100111000110000100101001110001101010011101101011010011"),
                ("10011100111101011010010011100010110101101101001001010011100001001010010100111000010010100101001010000100001000010000100001001010010100001001010011100011000100111001110011110101001110011100111001110110"),
                ("10011100111101011010010011100010110101101101001001010011100001001010010100111000010010100101001010000100001000010000100001001010010100001001010011100011000100111001110011110101001110011100111001110110"),
                ("10110100111001110011100111001110110101101001101001010011101001001010010100111000010010100001000010000100001000010000100001001010000100001001010010100111000100111011010110101101011010110101101011010110"),
                ("10011110011011010110101101011010110101101001111000110001001110110101101100001001010011100011000010010100001000010000100001000010011100011000110001101010011100111011010110101101011010110100111001110011"),
                ("11001110011011010110100111011010110101101011011010100111001110011100111101001001010011100011000010010100001000010010100101001010010100001001010011100011000100111011010110100111100111001110011100111001"),
                ("11001110011100111001110011001110110101101001110011101101101001001010011100001001010010100101001010000100001000010010100101000010000100001001010011100001001110101011010110110011100111001110011100101100"),
                ("11001110011100111001110011001110110101101001110011101101101001001010011100001001010010100101001010000100001000010010100101000010000100001001010011100001001110101011010110110011100111001110011100101100"),
                ("11001110011100111001110011100110110101101011010110110000100101001010011100001001010000100001000010000100001000010000100001000010000100001001010011100001001110101011010110110011100111001111011110101110"),

                -- explosion_1-1.png
                ("11111111111111011110011001100110011100111001110011101101001111000110000100111000100111001110011110101101011010010010100101001010011101011001110011100111001110011100111001110011100101100111111111111111"),
                ("11111111111100111001110011001110110101101011010110101101001101001010010100101001110101001110011010010100101001010000100001000010010100111010110101011010011100111001110011110011100111001111111111111111"),
                ("11111111111100111001110011100111001110011001110110101101101001001010011100001000010000100001000010000100101000010000100001000010011100011000110001101010011101101011010110110011100111001111111111111111"),
                ("11111111111100111001110011100111001110011001110110101101101001001010011100001000010000100001000010000100101000010000100001000010011100011000110001101010011101101011010110110011100111001111111111111111"),
                ("11111111110110001100011001100111001110011100110110101101001101001010010100101000010000100001000010010100001000010000100001000010011100010011100111001111010100111001110011110011100111001111111111111111"),
                ("11111111111111111111110011100111001110011100110110101101011010011100110100101000010000100101001010010100101001010010100101001010001100010011100111001111010100111001110011110011100111001111111111111111"),
                ("11111111111111111111111010110011001110011001110110101101001111010110100100101000010000100001000010010100101001010000100001000010001101010011100111101011010110011100111001110011100101100111111111111111"),
                ("11111111111111111111111010110011001110011001110110101101001111010110100100101000010000100001000010010100101001010000100001000010001101010011100111101011010110011100111001110011100101100111111111111111"),
                ("11111111111111011110111100110001100011001001110011110100100101001010010100101001010000100001000010000100001000010000100001001010011101011010110101100011010101101100111001110010110001100111111111111111"),
                ("11111111110111001110011001001111001110011001111000010010100111000110000100101001010010100101001010000100001001110101101011000010011101010011100111101011010101101011010110110011110101110111111111111111"),
                ("11111111111111111111011001011010110101101001101001010010100111000110000100101000010000100001000010000100001001110001100001001010011101011010110101101010011100111001110011110010110011111111111111111111"),
                ("11111111111111111111011001001110110101101011011000010011100011000110000100101000010000100001000010000100111000010010100101001010010100101001010011101010011101101011010110101101100111111111111111111111"),
                ("11111111110111001110011001100110110101101011011010010011101011000110000100101001010000100001000010010100101001010010100101001010010100101001010010100111010101101011010110101101001111001111111111111111"),
                ("11111111110111001110011001100110110101101011011010010011101011000110000100101001010000100001000010010100101001010010100101001010010100101001010010100111010101101011010110101101001111001111111111111111"),
                ("11111111111110111101110011100110011100111001111010110101001111010110100100101001010000100001000010000100101001010010100101001010010100111000110001001110110101101001110011100111001111001111111111111111"),
                ("11111111111100111001110011011010011100111101010011101101011011010110100100001000010000100001000010000100101001010010100111000110000100111010110101001111010100111001110011110011100111001111111111111111"),
                ("11111111111111011110111101100110110101101011010011100111001111010110100100101000010000100001000010000100001001010010100111010110000100101001010010100101001100111011010110101101100111101111111111111111"),
                ("11111111111111011110111101100111001110011011010110100111001111010110101101011000010010100001000010000100001000010000100001001010010100101001010010100111000101101011010110100111100101100111111111111111"),
                ("11111111111111011110111101100111001110011011010110100111001111010110101101011000010010100001000010000100001000010000100001001010010100101001010010100111000101101011010110100111100101100111111111111111"),
                ("11111111111110111101011001100110011100111100110110100111101011010110101100001001010010100001000010000100001000010010100101001010010100101001010010100111000100111100111001110011100101100111111111111111"),
                ("11111111110111001110011001100110011100111011010110101101011010011100111100001001010000100001000010000100001000010000100001001110000100101001010011101011000100111011010110110011100111001111111111111111"),
                ("11111111111110111101110011100111001110011100110011100111001110110101101101001001010010100001000010000100001000010000100001001010010100101001010011001110011100111011010110101101100111001111111111111111"),
                ("11111111110110001100110011100111001110011100110011110101001110011100111101001001010010100001000010010100001000010010100101001010010100101001010011001110110101101001110011101101100111001111111111111111"),
                ("11111111110110001100110011100111001110011100110011110101001110011100111101001001010010100001000010010100001000010010100101001010010100101001010011001110110101101001110011101101100111001111111111111111"),
                ("11111111111100111001110010110011001110011001110110100111101011010110100100111000010010100001000010000100001000010000100001000010010100101001010011101010011100111001110011101101001111001111111111111111"),
                ("11111111111111111111011000110010011100111011010110100111101001001010010100111000010000100001000010000100001000010000100001000010011101011010110101101011000110101011010110101101001111001111111111111111"),
                ("11111111111111111111111011100110110101101001110011100110100101001010011100001001010010100001000010000100001000110001100001001110001101011010110101001111000110101011010110101101001111001111111111111111"),
                ("11111111111111011110111100110011001110011001111000010010100111000110000100101001110100100101001010000100001000110001100001001010011101010011100111101010011110011100111001110011100111001111111111111111"),
                ("11111111111111011110111100110011001110011001111000010010100111000110000100101001110100100101001010000100001000110001100001001010011101010011100111101010011110011100111001110011100111001111111111111111"),
                ("11111111110110001100011001111001100011001011011010010010100101001010010100101001010010100101001010000100001000010010100101001010010100101001010011101010110110011100111001110011100111001111111111111111"),
                ("11111111111111111111011100110011001110011001111010100111101001001010010100001000010000100001000010000100001000010010100111000010010100101001010011101010110101101100111001110011100111111111111111111111"),
                ("11111111111111111111011100110011001110011001101001100111011011010110100100101001010000100001000010010100101000010010100111000010011001110011100111001110110100111100111001110010110011111111111111111111"),
                ("11111111111001110011011100110010011100111011001001110101011010011100110100101001010000100001000010010100101001110001100001001110001011010011100111101010110101101100111001011000111011110111111111111111"),
                ("11111111111001110011011100110010011100111011001001110101011010011100110100101001010000100001000010010100101001110001100001001110001011010011100111101010110101101100111001011000111011110111111111111111"),
                ("11111111110110001100011001100110110101101001101001100111011010011100111101001001010000100001000010000100001000010010100101001110001101011000110001100010011101101011010110110010110001100111111111111111"),
                ("11111111111110111101110011011010011100111001110110101101001111000110001101001000010000100001000010000100001000010000100001000010011100001001010011101010011110011001110011101101100111001111111111111111"),
                ("11111111111100111001100111011010110101101011010011100111101001001010010100101001010000100001000010000100001000010000100001000010010100101001010011100010011110011100111001110011100111001111111111111111"),
                ("11111111111100111001100111100111001110011001110011110100100101001010010100001001010000100001000010000100001000010000100001001010011100001001010011101010110101101011010110100111100101100111111111111111"),
                ("11111111111100111001100111100111001110011001110011110100100101001010010100001001010000100001000010000100001000010000100001001010011100001001010011101010110101101011010110100111100101100111111111111111"),
                ("11110011001100111001110011100110011100111100011000010010100101000010000100001000010000100001000010000100001000010010100101001110000100101001010011001110110101101011010110101101001101100111111111111111"),

                -- explosion_1-2.png
                ("11110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("01100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11001110011100111001111010110010011100111111111111011001111011111111111111111001011001110111101011101110111110111101111011001111010111011111111111111101110111101111111111111110110011001110011100111110"),
                ("11001110011100111001111010110010011100111111111111011001111011111111111111111001011001110111101011101110111110111101111011001111010111011111111111111101110111101111111111111110110011001110011100111110"),
                ("11001100111001110011110010110001110011100111001110011001111011101111010110011001110011100111001011000110011110111101111011001110010110001100011000110001100111101110111101110010110011001110011100101100"),
                ("11001110011011010110101101100101100011000110001100111100110011001110010110001100110011100111001110011100111001110011100110110110011100110011100111011010011011000110001100110011100111001100111001111001"),
                ("10011110011011010110100111011010011100111100111001011001100110110101101001111001110011100111001100111001111001101101011010011100111011010110101101011011001011001100111001110011100111001101101011010011"),
                ("10011110011011010110100111011010011100111100111001011001100110110101101001111001110011100111001100111001111001101101011010011100111011010110101101011011001011001100111001110011100111001101101011010011"),
                ("11000100111011010110100111001110110101101001110011101101001110011100111011010011110011100111001101101100110110101101011011010100111011010110101101001110011100111001110011110011100110011101101011010011"),
                ("11000100111001110011101100100101001010010100111010110101100010011100111011010110100111001110011101101011010110100111001110011110101101011000110000100111000100111011010110101101011010110101101011010011"),
                ("01001110101001110011101101001111010110101001110011010010100110011100111001110011110101001110011101101001110011100111001110110110100100101001010010100101001110101011010110101101011010110101101011010110"),
                ("01001010011101011010100111011010110101101011011010010010100101001010011101011010100111001110011101101101010011100111001110110100111101011000110000100101001010011001110011101101001111010100111001110011"),
                ("01000010010100101001110001001110011100111101001001010011100001001010010100111010100111011010110100111101011010110101101011010110101100011000110001100011000010011101011010100110100101001010010100111000"),
                ("01000010010100101001110001001110011100111101001001010011100001001010010100111010100111011010110100111101011010110101101011010110101100011000110001100011000010011101011010100110100101001010010100111000"),
                ("01000010000100101001110101101001001010010100101000010010100111000110000100101001110101101011010110001100011010010010100101000010010100101001010010100101001010010100101001010010100111000010010100101001"),
                ("01000010010100101001010000100101001010010100101000010010100101001010011100011000010010100101001010010100111000010000100001000010010100101000010000100001001010010100001000010000100001000010010100111000"),
                ("01000010000100001000010000100001000010000100001000010011101001001010010100001001010010100101001010000100101001010000100001000010000100001000010000100001001010000100001000010000100001000110101101010011"),
                ("01000010000100001000010000100001000010000100001000010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010000100001000010010100001000100111001110011"),
                ("01000010000100001000010000100001000010000100001000010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010000100001000010010100001000100111001110011"),
                ("01000010000100001000010000100001001010010100101000010000100001000010000100001000010010100001000010000100001000010000100001000010000100101000010000100001000010000100101001010010100101000010010100111010"),
                ("01000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001010010100001000010000100101001010010100001001010010100111010"),
                ("01000010000100001000010000100001001010010100001000010000100001000010000100001000010000100001000010000100001000010010100101001010010100111000110000100101001010000100101001010010100001000010010100111010"),
                ("01001010000100001000010000100111000110000100101001010011100011000110000100001000010010100001000010000100101000010010100101001010010100101001010011100011010010000100001000010010100001000010000100001001"),
                ("01001010000100001000010000100111000110000100101001010011100011000110000100001000010010100001000010000100101000010010100101001010010100101001010011100011010010000100001000010010100001000010000100001001"),
                ("01001010010100001000010000100101001010011100011000010010100101001010010100001000010010100101001010010100101001110101101011000010010100101001010010100111000010010100001000010010100001000010000100001001"),
                ("11000010010100101001010011100011000110000100101001010010100111000110000100101001010010100101001110000100101001110001100011000010010100101001010010100101001010010100001000010000100101001010010100101001"),
                ("01001110000100101001110001101010110101101001101001010011101011010110101101001001010010100101001010010100101001010010100101001010010100101001010011101011010110101101011010110001100011000010010100111010"),
                ("01001010010100101001010011100010011100111001101001010011001111010110101101001001010010100101001010010100101001010010100111010110000100101001010011101010011110101001110011100111001111000110101101011001"),
                ("01001010010100101001010011100010011100111001101001010011001111010110101101001001010010100101001010010100101001010010100111010110000100101001010011101010011110101001110011100111001111000110101101011001"),
                ("10011110101100011000110101100011010110101001111010110101101010011100111101011010100111001110011110100100101001010010100110011100110100111010110101101011010110001101011010100111001111010101101011011001"),
                ("10110101101001110011100111001110110101101011010110101101001111000110001100010011101101001110011110001100011000010010100111010101101101010011100111001111010110101101011010110101101010011100111001111001"),
                ("10110101101100111001110011011010110101101001110110110011100111010110101101010011101101001110011100111001110110100111001110011101101011010110101101001110110101101100111001100111001110110100111001111001"),
                ("10110101101100111001100111011011001110011100111001110011100110110101101011010011100111011010110101101100110110101101011010011100111011010110101101001110110110011100111001100111001110110100111001111001"),
                ("10110101101100111001100111011011001110011100111001110011100110110101101011010011100111011010110101101100110110101101011010011100111011010110101101001110110110011100111001100111001110110100111001111001"),
                ("10110100111100111001101101100101100011001100111001110011100110110101101011010110101101011010110110011100110011101101011011001100111011010110101101100111001110011100111001110011100111001110011100111001"),
                ("10011110011100111001110010110001110011100110011001110011100110011100111001110011110011100111001110011100111001110011100111001100111001111001110010110011101011001100111001110011100111001110011100111001"),
                ("01100011001100111001110010110011110111101111111111110011100111001110011100111001110011100111001110010110001100111011110111001110011100111111111111111101110011000110001100110011100111001110011100101100"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_1-3.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010110101101010011110101001110011100111001111001111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111001100111001110011110010110001100111101111011001111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111100111001101101011010110100111100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111100111001101101011010110100111100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111110111101100111001110011001110011101101011010110101101011011001110011100111001110011100101100011000111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111101100111101100111001110011011010110101101011010110101101011010011100111001111001110011100111001110010110011101111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111110101100110011100111001110011001110011100111011010110100111001110110101101011010110110011100111001110011100101100111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111110101100110011100111001110011001110011100111011010110100111001110110101101011010110110011100111001110011100101100111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111001110011100101100110011100111001110011001110011101101011010110101101001110110101101011010110101101100111001110011100111001110011001110011111111111111111111111111111111"),
                ("11111111111111111111111110110010011100111011011001110011100110011100111011011010100111011010110101101011010110101101011010110101101100110011100111011010110101101001110011011001111111111111111111111111"),
                ("11111111111111111111111111100111001110011011010011101101011010011100111001111010110101011010110101101001110011100111001110011100111001110011100111011010110101101001110011110011110111111111111111111111"),
                ("11111111111111111111111111100111001110011001110110101101011011010110101101011000110101001110011100111001101001110101101011000010011100010011100111011010110100111100111001110010110011110111111111111111"),
                ("11111111111111111111110011100110011100111001110110101101001101001010010100111010110101101011010100111101001001010010100101001110101101011010110101001110110101101001110011110011100101100111111111111111"),
                ("11111111111111111111110011100110011100111001110110101101001101001010010100111010110101101011010100111101001001010010100101001110101101011010110101001110110101101001110011110011100101100111111111111111"),
                ("11111111110110001100110011011010011100111100110011101101101001001010010100111000100111001110011110100100101001010010100111010101101001111000110001101010110101101001110011110011100111111111111111111111"),
                ("11111111111100111001110011011010011100111100111001101101001111010110101101001001110101100011000010010100101001110101101011010101101001111000110001101010110101101001110011101101011011111111111111111111"),
                ("11111111111100111001110011100110011100111001110011110101101011010110101100001001010010100101001010000100101001110001100011000110100100101001010011101010110101101011010110101101001111001111111111111111"),
                ("11111111111100111001110011100110011100111011010011010010100111010110100100111000010010100101001010000100111000010010100101001010011101011000110001001110110101101011010110101101100111001111111111111111"),
                ("11111111111100111001110011100110011100111011010011010010100111010110100100111000010010100101001010000100111000010010100101001010011101011000110001001110110101101011010110101101100111001111111111111111"),
                ("11111111111100111001110011001110110101101001110011110000100101001010010100101001110000100101001010000100001001010010100101001110001001110110101101011010110101101011010110100111100111001111111111111111"),
                ("11111111111100111001110011011010110101101011010011110000100101001010010100111000010010100101001010000100001000010010100111000010011101010110101101001110110101101001110011110011100111001111111111111111"),
                ("11111111111100111001110011100110110101101011010110110100100101001010010100101001010000100001000010000100001000010010100111000010010100111010110101100011010101101011010110110011100111001111111111111111"),
                ("11111111111100111001110011001110011100111101011010100111101010011100111101001001010000100001000010000100001000010010100111000010011100011010110101101001001100111011010110110010110001100111111111111111"),
                ("11111111111100111001110011001110011100111101011010100111101010011100111101001001010000100001000010000100001000010010100111000010011100011010110101101001001100111011010110110010110001100111111111111111"),
                ("11111111111100111001110011011011010110101001110110101101011010110101101101001001010011100011000010000100001000010010100111000010011001110110101101001111010110101011010110110011110111111111111111111111"),
                ("11111111111100111001110011001111010110101101010011100111101011000110000100101001010010100101001010000100001000010010100111000010011101010011100111001110110100111011010110100111100111111111111111111111"),
                ("11111111111100111001110011001111000110001100010011110100100101001010010100111000010010100001000010000100001001010010100101001010010100111000110001101010110101101011010110100111100101100111111111111111"),
                ("11111111111100111001110011001110011100111001110011010010100101001010010100111000010010100101001010000100001001010000100001000110000100111010110101001110110101101001110011110011100111001111111111111111"),
                ("11111111111100111001110011001110011100111001110011010010100101001010010100111000010010100101001010000100001001010000100001000110000100111010110101001110110101101001110011110011100111001111111111111111"),
                ("11111111111111111111110011100110011100111011010011010010100101001010010100101001010010100101001010000100001000010000100001000010011100011010110101001111001110011100111001110011100111111111111111111111"),
                ("11111111111111111111011001100111001110011001110110100111101001001010010100101001010000100001000010000100001000010000100001001110001100010011100111001110011110010110001100011001100111111111111111111111"),
                ("11111111110110001100110011100110011100111011010110101101011011010110100100111000010010100001000010000100001000010010100101001010011100010011100111101010110100111100111001011001100111001111111111111111"),
                ("11111111111100111001110011100110011100111011010110101101001111010110100100101001010000100001000010000100001000010010100101001010011101010110101101001111010100111100111001110010110001100111111111111111"),
                ("11111111111100111001110011100110011100111011010110101101001111010110100100101001010000100001000010000100001000010010100101001010011101010110101101001111010100111100111001110010110001100111111111111111"),
                ("11111111111100111001110011001110110101101011010110101101001111000110000100101001010000100001000010000100001000010010100101001010011001110110101101001101001110101100111001011001111001100111111111111111"),
                ("11111111111100111001110011100110110101101011010110101101011011010110100100101000010000100001000010000100001000010010100101001010011001110110101101011010011100111001110011011001111011101111111111111111"),
                ("11111111111100111001110011100110011100111011010110101101011010011100110100101001010010100001000010000100001000010000100001001010011101010110101101011011010010011001110011110010111011110111111111111111"),
                ("11111111111100111001110011100111001110011011010110101101011010110101101101001001010000100001000010000100001000010000100001001010011101010110101101011010011110101001110011110010110001100111111111111111"),
                ("11111111111100111001110011100111001110011011010110101101011010110101101101001001010000100001000010000100001000010000100001001010011101010110101101011010011110101001110011110010110001100111111111111111"),
                ("11111111111111111111110010110001100011001100110110101101011010011100111101001001010010100101001010010100001000010000100001000010011001110110101101011010011101101100111001011001111111111111111111111111"),

                -- explosion_1-4.png
                ("11111111111111111111111110110011001110011011010011101101011010011100110100101000010000100001000010000100101001010010100101001110101001110110101101011010110110010110001100011001100111111111111111111111"),
                ("11111111110110001100011001100110011100111101010011101101011011010110100100101001010000100001000010000100001000010000100001001110101011010110101101011010110101101100111001110011100111001111111111111111"),
                ("11111111111111011110011101100110011100110100111010101101011011010110100100101001010000100001000010000100001000010010100101001010011001110110101101011010110101101001110011110011100111001111111111111111"),
                ("11111111111111011110011101100110011100110100111010101101011011010110100100101001010000100001000010000100001000010010100101001010011001110110101101011010110101101001110011110011100111001111111111111111"),
                ("11111111111110111101111100110010011100111001110011101101011010011100110100101001010010100001000010000100001000010000100001000010011101010110101101011010110101101011010110110011100111001111111111111111"),
                ("11111111110110001100111100110011001110011101001001100111011010011100110100101001010010100001000010000100001000010000100001001010011100010011100111011010110101101011010110100111100111001111111111111111"),
                ("11111111110110001100011001100111001110011001111010100111011011010110100100101001010010100001000010000100001000010000100001001010011101010011100111011010110101101001110011110011100111001111111111111111"),
                ("11111111110110001100011001100111001110011001111010100111011011010110100100101001010010100001000010000100001000010000100001001010011101010011100111011010110101101001110011110011100111001111111111111111"),
                ("11111111111100111001110010110011001110011001110110110101001111000110000100101001010010100001000010000100001000010010100111000010011101010110101101011010110101101001110011110011100101100111111111111111"),
                ("11111111111111111111110010110001100011001100110011100111001111000110001100001001010000100001000010000100001000010000100001001010010100111010110101001110110100111100111001110010110011111111111111111111"),
                ("11111111111111111111110011100111001110011100111001100111101011000110000100101000010000100001000010000100001001010010100101001010010100101001010010100110011101101001110011110011100111111111111111111111"),
                ("11111111111100111001110011100110011100111011010110100111101001001010011100001000010000100101001010000100001001010010100111000010010100101001010010100110011100111001110011100111100111001111111111111111"),
                ("11111111110110001100110011001110110101101011010110110101100001001010010100101001010010100101001010000100001000010010100111000010010100101001010011101010011110001100011000100111100111001111111111111111"),
                ("11111111110110001100110011001110110101101011010110110101100001001010010100101001010010100101001010000100001000010010100111000010010100101001010011101010011110001100011000100111100111001111111111111111"),
                ("11111111111111111111110011001110110101101001110110100111001111010110100100111000010010100001000010000100001001010010100101001010011100011010110101001110011110101101011010100111100111001111111111111111"),
                ("11111111111111111111111011100110110101101101011010100111011010011100110100111000010010100001000010000100011000010010100101001110101011010110101101011010110100111101011010101101100111001111111111111111"),
                ("11111111110110001100011001100110110101101001101001110101101011000110000100111000010010100001000010000100001000010000100001001110101001111010110101001111010110101001110011100111100111001111111111111111"),
                ("11111111111100111001110011100110110101101011011010110001101001001010010100111000010010100001000010000100001000010000100001001010010100101001010011101010110101101011010110110011100111001111111111111111"),
                ("11111111111100111001110011100110110101101011011010110001101001001010010100111000010010100001000010000100001000010000100001001010010100101001010011101010110101101011010110110011100111001111111111111111"),
                ("11111111111100111001110011100110011100111011010110100111011011010110100100111000010010100001000010000100001001010010100111000010010100101001010011100010011101101011010110101101100111001111111111111111"),
                ("11111111111100111001110011001110110101101011010110101101011010011100111100001001010010100101001010000100001001110001100001001010010100101001010011100010011100111011010110100111100111001111111111111111"),
                ("11111111111100111001110011011010110101101011010110100111100011010110100100101001010011100011000010010100001001010010100111000010011101001001010010100110011101101001110011110011100111001111111111111111"),
                ("11111111111100111001100111011010110101101011010110110100100101001010011101011000110000100101001010010100001001010010100101001110001101011010110101101010011100111001110011110011100111001111111111111111"),
                ("11111111111100111001100111011010110101101011010110110100100101001010011101011000110000100101001010010100001001010010100101001110001101011010110101101010011100111001110011110011100111001111111111111111"),
                ("11111111111111111111101101011010011100111011010110110101100010011100111011011010110100100101001010010100111000110101101001001110101101010011100111011011001110011001110011101101100111001111111111111111"),
                ("11111111111111111111110011100110011100111011010110110101100010011100111011011010010010100101001010011101010011100111001111000010010100111010110101011010011110011001110011101101100101100111111111111111"),
                ("11111111110110001100110011100110011100111011010110100111101011010110101101001001010010100101001110101001111010110101101011010010010100110011100111011010110100111001110011110011100111111111111111111111"),
                ("11111111111111011110011001100111001110011001110110101101001111000110000100111000110100100101001100111001110011110101101011000110101101010110101101011010110100111100111001110011111111111111111111111111"),
                ("11111111111111011110011001100111001110011001110110101101001111000110000100111000110100100101001100111001110011110101101011000110101101010110101101011010110100111100111001110011111111111111111111111111"),
                ("11111111111111111111111011100110011100111011010110101101001110011100111001110011100111001110011100111011010110110101101011010100111001110110101101011010011101101100111001110011111111111111111111111111"),
                ("11111111111111111111111110110010011100111011010110101101001111001110011011010110101101011010110101101011010110100111001111010101101001111001110011100111001101101001110011011001111111111111111111111111"),
                ("11111111111111111111111111111110011100111100111001110011100111001110011011010110101101011010110100111011010110101101011010011100111100111001110011100101100110011100111001111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111001100110011100111001110011100110110101101011010110100111001110110100111001110011100111100111001110011100101100111011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111001100110011100111001110011100110110101101011010110100111001110110100111001110011100111100111001110011100101100111011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111101011001100111001110011100111001100111001110011101101011010110101101011010110101101100111001110011111001100111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111011100110011001110011100111001110011100111001101101011010110101101011010011100111100111001110011111011110111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111100111001110011100111001110011001110110101101011011001110011111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111001111100110001100011001100110011100111001111001111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111001111100110001100011001100110011100111001111001111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111001100111001110011100111101010011110101101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_1-5.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111110011100111001110011100111001110010110011111111111100111001110011100111001110011100111001110011100111001110011100111001011001111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111110011100111001110011100111001110010110011111111111100111001110011100111001110011100111001110011100111001110011100111001011001111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11001110011100111001110011100111001110011100101100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111"),
                ("01100110011100111001110011001111001110011100111001110011001110011100111001110110100111100111001101101001111001110011100110110101101100111001110011100101100111111111111111111111111111111111111111111111"),
                ("01100110011001110011101101011010011100111001111001100111001111000110001101011010100111011010110101101011010011100111001110011100111001111001110011100110011110011111111111111111111111111111111111111111"),
                ("01100110011001110011101101011010011100111001111001100111001111000110001101011010100111011010110101101011010011100111001110011100111001111001110011100110011110011111111111111111111111111111111111111111"),
                ("11001101101011010110101101011010110101101011010011101101001111000110001101010011110101011010110101101001110110100111001111001110011001110011100111011010110110011110111101111111111111111111111111111111"),
                ("10110101101011010110101101011010110101101011010110100111001110011100111001110110110101011010110100111001110011100111001111001100111011010110101101001111001011000110001100011001111011111111111111111111"),
                ("10110101101011010110101101011010110101101011010011010010100111010110101001110110100111101011010110001100001001110101101010110101101011010110101101011011001110011100111001111101111011111111111111111111"),
                ("10110101101011010110101101001110011100111011011010010010100101001010011101010110110100100101001010010100101001110101101010011110101001110110101101011011001110011100111001110011100111111111111111111111"),
                ("10011101101001110011110101100011010110101101001001010010100101001010011100010110100110100101001010010100111010110101101011010010010100111010110101001110011110011100111001110011100111111111111111111111"),
                ("10011101101001110011110101100011010110101101001001010010100101001010011100010110100110100101001010010100111010110101101011010010010100111010110101001110011110011100111001110011100111111111111111111111"),
                ("11010110100100101001010010100101001010010100101001010010100101001010010100111010110100100101001010010100101001110001100011010010010100111010110101001110110100111001110011101101001111001111111111111111"),
                ("01001010010100101001010000100101001010011100001001010011100011000110000100101001010010100101001110000100111000010010100101001110001101011000110001101011010100111001110011101101001111001110011100111111"),
                ("01001010000100101001010000100001000010000100101000010010100101001010010100101001010000100001000010011100001001010010100111010100111101011010110101101010011101101001110011101101011010110100111001111111"),
                ("01001010000100001000010000100001000010000100001000010010100101000010000100111000010000100001000010010100101001010010100111000100111101010011100111011010110101101011010110101101011010110100111001111111"),
                ("01001010000100001000010000100001000010000100001000010010100101000010000100111000010000100001000010010100101001010010100111000100111101010011100111011010110101101011010110101101011010110100111001111111"),
                ("01001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001110101001110011100111011010110101101001110011101101011010011110011100111111"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001010011101010011100111001110110100111001110011101101011011001011000110011111"),
                ("01000010000100001000010000100001000010000100001000010000100101001010010100001000010000100001000010000100111000010010100101001010010100101001010011001110110101101011010110100111100111001011000110011010"),
                ("01000010000100001000010010100101001010010100101000010000100001001010010100101001010010100101001010010100101001110001100011010010010100111010110101001110110101101011010110100111100111001111101111011010"),
                ("01000010000100001000010010100101001010010100101000010000100001001010010100101001010010100101001010010100101001110001100011010010010100111010110101001110110101101011010110100111100111001111101111011010"),
                ("01000010010100101001010010100101001010010100101001010000100001001010011100011000110001100011000110000100101001110001100011010110100100111000110001001110110101101011010110110011100111001110011100110011"),
                ("01001010010100101001010010100101001010010100111000010011100001001010010100101001010010100101001010011100001001110101101010110101101101001001010011001110110101101100111001110011100111001111111111111010"),
                ("10011110101101011010100111001111010110101100011000110000100101001010011101010011110000100101001110101001111010010010100110011100111101011000110001001111001110011100111001110011100111111111111111110011"),
                ("10110101101011010110101101011010110101101001110011110101101011000110001001110110110101101011010101101011011000010010100111000110001101010011100111001110011110011100111001110010110011111111111111110011"),
                ("10110101101011010110101101011010110101101001110011110101101011000110001001110110110101101011010101101011011000010010100111000110001101010011100111001110011110011100111001110010110011111111111111110011"),
                ("10110101101011010110101101001110011100111101010011100111001111010110101001110011110101100011000100111011010011110101101011010110101001110110101101011010110110011100111001011000111011111111111111110011"),
                ("10011100111101011010100110100111010110101011010011110011011010110101101011011010010011101011010101101011010110101101011010110101101011010110101101011010110110010110001100111011111111111111111111111001"),
                ("10110110100100101001100111101010011100111001111001110011011010110101101001111010100111011010110101101011010110101101011010110101101011010011100111011010110110011111011110111111111111111111111111111111"),
                ("11001100111001110011100111100111001110011100101100110011001110110101101011010110101101011010110100111011010110101101011010011100111001111001110011001110011100111111111111111111111111111111111111111111"),
                ("11001100111001110011100111100111001110011100101100110011001110110101101011010110101101011010110100111011010110101101011010011100111001111001110011001110011100111111111111111111111111111111111111111111"),
                ("01100110011100111001011000110011001110010110001100110011100110011100111001111001110011100111001110011001110110101101011010110110011100111001110011100101100111111111111111111111111111111111111111111111"),
                ("11111011000111001110111101111001100011001100111001110011100111001110011100111101011001100111001110011100111001100111001110110110011100101100011001110111111111111111111111111111111111111111111111111111"),
                ("11111011001111011110111010110001100011001100111111111111100101100011001111111111011001100111001110011100111001110011100111111111110110011110111101111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_1-6.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111001100011001111111111110011100111001110011100111001011000110011111111110110011001110011111111111110010110001100011001110111110011000110011111"),
                ("11111111111111111111111111111111111111111111111111111111111001100011001111111111110011100111001110011100111001011000110011111111110110011001110011111111111110010110001100011001110111110011000110011111"),
                ("11111111111111111111111111111111111111111111111111111010110011001110011100110110100111100111001110011100111001011000110011101110011100111001110011100111001110010110001100111101111001110011000110011111"),
                ("11111111111111111111111111111111111111111111101100110011100111001110011100110110101101011010110100111100111001110011100111001100111001111001110011100101100011001100111001011000110011001110011100101100"),
                ("11111111111111111111111111111111111111111001110011100111100110011100111001110011101101011010110101101001110110101101011010110101101011010011100111100101100110011100111001110011001110011100111001111001"),
                ("11111111111111111111111111111111111111111001110011100111100110011100111001110011101101011010110101101001110110101101011010110101101011010011100111100101100110011100111001110011001110011100111001111001"),
                ("11111111111111111111111111111111110111101100110110101101001110110101101011010110101101011010110101101011010110100111001111010100111011010110101101100111001100111001110011110101001101001110101101010110"),
                ("11001111111111111111111111110101100011001100110110101101011010110101101011010110101101011010110101101011011010010010100111010101101011010110101101100110011101101101011010010011001111010100111001110011"),
                ("10011111111111111111011100110011001110011100110110101101011010011100111101011010110101001110011101101001111000110101101010011100111101010011100111001110011110101001110011100111011010110101101011010110"),
                ("10011111111111111111011001100111001110011100110011100111001111010110101100011000010011100011000101101011011010110101101010110100111100011010110101101010011100111011010110101101011010110101101011010110"),
                ("10011111111111111111110011100111001110011100111001100111100011010110101001110011010011101011010100111101001001110001100010011110100100101001010011100011000110001101011010100111001111010110101101010011"),
                ("10011111111111111111110011100111001110011100111001100111100011010110101001110011010011101011010100111101001001110001100010011110100100101001010011100011000110001101011010100111001111010110101101010011"),
                ("11010111111100111001110011100111001110011011010110100110100111010110101011010110110100100101001110000100101001010010100101001010010100111000110000100111000010010100101001010010100101001010010100101001"),
                ("10011110011100111001110011100110110101101011010110100111100001001010011101011010110000100101001010011100011000110001100011000110000100101000010000100001001010010100101001010010100101001010010100101000"),
                ("11010111101100111001110011001110110101101011010110100111101001001010010100111010110000100101001010010100101001010010100101001010010100101000010000100001000010010100101001010010100101000010000100001000"),
                ("11010011001100111001110011001110110101101011010110100110100101001010010100101001010011100011000010010100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001000"),
                ("11010011001100111001110011001110110101101011010110100110100101001010010100101001010011100011000010010100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001000"),
                ("11111011001100111001101101011010011100111001110110100111001111010110100100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("11111110011001110011101101011010011100111011010110101101001110011100111101001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001"),
                ("11111100111011010110101101011010110101101011010110101101001111010110101001111000010010100101001010010100101000010000100011000010010100001001010010100101000010000100001000010000100001000010000100001001"),
                ("11111100111011010110101101011010011100111011010011110101101011010110101001111010010010100101001110000100101000010000100001001010010100101001010010100101000010010100001000010000100001001010000100001001"),
                ("11111100111011010110101101011010011100111011010011110101101011010110101001111010010010100101001110000100101000010000100001001010010100101001010010100101000010010100001000010000100001001010000100001001"),
                ("11111110011100111001100111011010011100111001111010110101100011010110101100001001010011100011000010011100001001010010100101001010011100011000110000100101001110000100101001010010100001001010010100101001"),
                ("11111111111100111001100111011010011100111001110110100111101001001010010100111010110000100101001010010100101001110101101011010010010100101001010010100101001010010100101001010010100101001110101101011010"),
                ("11111111111111111111110011100111001110011100110011100111101001001010010100111010110101101011010010010100101001100111001110110110000100101001010010100101001110101101011010110001101010011101101011010011"),
                ("11111111111111111111110011100111001110011100111001101101011010011100111101010011110100100101001010010100101001110101101010110110100100101001010010100111010101101001110011100111011010110101101011010110"),
                ("11111111111111111111110011100111001110011100111001101101011010011100111101010011110100100101001010010100101001110101101010110110100100101001010010100111010101101001110011100111011010110101101011010110"),
                ("11111111111111111111111101111011001110011100111001101101011010110101101011010110110100100101001110001100011010100111001110110100111101001001010010100110011101101011010110101101011010110101101011010110"),
                ("11111111111111111111111100110001100011000110011001100111011010110101101001111001100111001110011100111001110110110101101010110100111001110011100111001110110101101011010110101101011010110101101011010110"),
                ("11111111111111111111111111111111101111011100110110101101001110011100111100111001100111011010110100111011010110110101101010011110101100010011100111011010011101101011010110101101011010110101101011011001"),
                ("11111111111111111111111111111111111111111100110011110011100110011100111001110011100111001110011101101011010110100111001111010110101100010011100111001111001100111001110011101101011010011110011100101100"),
                ("11111111111111111111111111111111111111111100110011110011100110011100111001110011100111001110011101101011010110100111001111010110101100010011100111001111001100111001110011101101011010011110011100101100"),
                ("11111111111111111111111111111111111111111111101100110011100111001110011011010110110011100111001100111011011001100111001110110100111001110011100111100111001110011100111001100111100111001110011100101100"),
                ("11111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100101100110011100111001110011100111001110011100111001"),
                ("11111111111111111111111111111111111111111111111111111111111111111111110110011001110011100111001110011100111001110011100111001110011100111001110011111111111011001100111001110011100111001110011100111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_2-0.png
                ("11111110010110001100110011100110110101101001111000010010100001000010000100001000010000100001000010001101111011010000100001000010000100111000110001101011000110101011010110011001111001100111101111011110"),
                ("11111110010110001100110011100110110101101101001000010000100001000010000100001000010000100001000010001011100001010000100001000010000100101001010010100110011100111011010110110010110011101110011100101100"),
                ("11001011000110001100110011100110011100111001101001010010100101000010000100001000010000100001000010001011100001010000100001000010000100111000110000100110011101101011010110100111100111001110011100111001"),
                ("11001011000110001100110011100110011100111001101001010010100101000010000100001000010000100001000010001011100001010000100001000010000100111000110000100110011101101011010110100111100111001110011100111001"),
                ("01100011001100111001110011100111000110001101011010010010100101000010000100001000010000100001000010001011100001110111101101000010000100001001010011100011000100111011010110101101100110011110011100111001"),
                ("10011110011100111001110011100111000110001101011010010010100001000010000100001000010000100001000010001101110111101111011110111010000100001001010010100101001110101001110011100111011010110101101011010011"),
                ("10110100111100111001110011101011010110101001111010010010100001000010000100001000010001011110111101111011101000010000100001000010000100001000010000100001000010011101011010101101011010011101101011001100"),
                ("10110100111100111001110011101011010110101001111010010010100001000010000100001000010001011110111101111011101000010000100001000010000100001000010000100001000010011101011010101101011010011101101011001100"),
                ("10110101101011010110100111101010011100111001111010010010100001000010000100001000101110000100001000010000111011010000100001000010010100101001010010100001000110001001110011110101101011000110101101001100"),
                ("10011100111101011010110101101010110101101101001001010000100001000010000100001000101110000100001000011011100001101111011101000010000100001000010000100101001110101101011010010010100001001010010100111000"),
                ("01001010010100001000010001100010011100111100001001010000100001000010000100001000101110000100001101110100011011101111011101000010000100001000010000100111010010010100101001010010100111000010010100101000"),
                ("01001010000100001000010000100111000110000100001000010000100001000010000100001000110111101111011010000100001000101111011101000010000100001000010001101011010110001100011000010011100011000110001100001000"),
                ("01000010000100001000010000100001001010010100001000010000100001000010000100001000010000100001000101111101110111101111011101000010000100001000010001100001001010010100101001010010100101001010010100101001"),
                ("01000010000100001000010000100001001010010100001000010000100001000010000100001000010000100001000101111101110111101111011101000010000100001000010001100001001010010100101001010010100101001010010100101001"),
                ("01000010000100101001010000100001000010000100001000010000100001000010000100001000010000000100001000011011101000110111101101000010000100001000010000100101000010000100001000010000100001000010000100001000"),
                ("01000010000100001000010010100101000010000100001000010000100001000010000100001000010001101111011000011011111011101111011111011010000100001001010010100001000010000100001000010000100001001110001100001000"),
                ("01000010000100001000010000100010111101111101101000010000100001000010000100001000010000100001000010000000110111101111011111011010000100001000010000100011011101110100001000010000100011000100111001101000"),
                ("01000010000100001000010001101100001000011101101000010000100001000010000100001000010001101111011101110000100001110111101101000010000100001000010000100011011110111101111011110111101101000010000100001000"),
                ("01000010000100001000010001101100001000011101101000010000100001000010000100001000010001101111011101110000100001110111101101000010000100001000010000100011011110111101111011110111101101000010000100001000"),
                ("01000010000100001000010001101111011110111011110111010000100001000010000100001000101111011110111000010000100001101111011101000010000100001000010000100001000101111011110111101111011101000010000100001000"),
                ("01000010000100001000010000100001000010001011110111101110100001000010000100011011101110100001000101110000100001000010000111011010000100001000010000100001000101111011110111000011011101000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000110111011110111110111011100001101111011100001010000100001000010000100001000010001101111011101111101101000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100000001101110100001000110111011110111010000100001000010000100001000010000100001000010001011110111101111101101000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100000001101110100001000110111011110111010000100001000010000100001000010000100001000010001011110111101111101101000010000100001000"),
                ("01000010010100101001010000100001000010000100001000010000100001001010011101100001010000100001000101111101110111010000100001000010000100001000010000100001000010000100001000010000100001001010000100001000"),
                ("01000010011101011010010010100001000010000100001000010010100101001010011101110111110111101111011110110100001000110111101101000010000100001000010000100001000010000100001000010000100001001010010100100011"),
                ("01001010011100011000010010100001000010000100001000010011101001001010010100011011000011011110111010001101110111010000100001000010000100001000010000100001000010000100001000010000100101001010000100011110"),
                ("01000010011100011000010010100101001010011100001001010000100101000010000100001000110111011110111101111011100001110111101101000010000100001000010000100001000010000100001000010000100101001110001100011110"),
                ("01000010011100011000010010100101001010011100001001010000100101000010000100001000110111011110111101111011100001110111101101000010000100001000010000100001000010000100001000010000100101001110001100011110"),
                ("01000010000100101001010010100101001010011001111010010000100001000010000100001000110110000100001000010000110111101111011101000010000100001000010000100001001010010100101001010000100001000110001100011110"),
                ("10011010010100001000010001100011010110101101001001010010100001000010000100001000110110000100001000010000101000010000100001000010000100001000010000100011000110001101011010110100100001001011000110001100"),
                ("10110110100100001000010001001110011100111101001000010010100101000010000100001000010001011110111110111101101000010000100001000010000100001000010000100111000010011101011010110101101011000110011100101100"),
                ("10110110100100001000010011011010110101101101001000010011101001001010010100001000010000100001000110110100001000010000100001000010000100111010110101001111010110101101011010110101001110110110011100111001"),
                ("10110110100100001000010011011010110101101101001000010011101001001010010100001000010000100001000110110100001000010000100001000010000100111010110101001111010110101101011010110101001110110110011100111001"),
                ("11001101101101011010100111011010011100111001101001010000100111000110000100101000010001011110111000010000111011010000100001000010000100011010110101001110011100111101011010110101001110110110011100111001"),
                ("10011101101011010110100111011010110101101001110011010000100101001010010100011011101110000100001000011011101000010000100001001010000100011000110001001110011100111100011000100111100110110110011100111101"),
                ("10110101101011010110101101011010110101101001110011110100100101000010001101100001000010000100001000010000101000010000100001001010010100001001010010100111010100111101011010100111100111001110011100111110"),
                ("11111100111100111001101101011010110101101011010011110100100101000010001011100001000010000100001110110100001000010000100001000010011100011000110000100111010101101001110011101101100101100011000110011110"),
                ("11111100111100111001101101011010110101101011010011110100100101000010001011100001000010000100001110110100001000010000100001000010011100011000110000100111010101101001110011101101100101100011000110011110"),
                ("11111111110110001100110011100111001110011011011010010010100001000010001011100001000010000100001101111011111011010000100001000010000100111000110000100111010101101011010110110010110001110111111111111111"),

                -- explosion_2-1.png
                ("11111011000110001100110011001110110101101001111000010010100001001010010100001000110111101111011101111101101000010000100001001010011101001001010010100111010100111011010110101101011011001111101111011111"),
                ("11111011001100111001110011001110110101101001111010100111100001001010010100001000010001101111011000011011101000010000100001001010011101001001010010100111010110101001110011101101011010011011000110011111"),
                ("11111110011100111001110011001110110101101011010011100111101001001010010100001000010000100001000101111011100001101111011101000010000100001000010000100111010100111001110011110101011011001110011100111111"),
                ("11111110011100111001110011001110110101101011010011100111101001001010010100001000010000100001000101111011100001101111011101000010000100001000010000100111010100111001110011110101011011001110011100111111"),
                ("11111011000110001100110011011010110101101011011010010011100001000010000100001000010001101111011101111011110111000010000110111010000100001000010000100001000010011100011000110101011011001011000110011111"),
                ("11111111101110111101011001011010110101101001111000010010100101000010000100001000010000100001000110111011100001110111101101000010000100001000010000100001000010010100101001100111011001100011100111011111"),
                ("11111111111111111111111101001110110101101011011010010010100101000010000100001000010000100001000101111011100001010000100001000010000100001000010000100111010100111011010110101101011001100011100111011111"),
                ("11111111111111111111111101001110110101101011011010010010100101000010000100001000010000100001000101111011100001010000100001000010000100001000010000100111010100111011010110101101011001100011100111011111"),
                ("11111111111111111111111101100110011100111011010110110100100001000010000100001000010000100001000010001101100001010000100001000010000100001000010000100001001110101011010110101101100101100111111111111111"),
                ("11111011001111011110111011100110110101101011010110100110100001000010000100101001010000100001000010000100010111110111101111011010000100001000010001101011010110101011010110101101100111110111111111111111"),
                ("11111010010110001100110011100110110101101011010011100111100001000010000100101000010001011110111110110100001000110111101110111010000100011000110001001110110100111011010110101100110011110110011100111111"),
                ("11111010001001110011110011011010110101101001111000010010100001000010000100101000010000000100001000010000100001000010000110111110110100001000010000100111010100111101011010100110110011001100111001111111"),
                ("11111010001100111001110011001110011100111001101001010010100001000010000100001000010000000100001000010000100001000010000100001101110100001000010000100001001110101001110011100111100111001110011100111111"),
                ("11111010001100111001110011001110011100111001101001010010100001000010000100001000010000000100001000010000100001000010000100001101110100001000010000100001001110101001110011100111100111001110011100111111"),
                ("11111010000001100011011000110011010110101001110011110100100111000110000100001000010001011110111101111011100001101111011110111110110100001001010010100001000100111011010110100110110011001011000110011111"),
                ("11111010001101011010110101100110011100111101010110100111101011000110000100101000110110000100001101110000100001110111101101000010000100001001010010100110011101101001110011110011100111001111101111011111"),
                ("11111110001100111001101101100110011100111011010110100110100101001010010100101000010001011110111000011011110111010000100001000010000100101000010000100110110101101011010110101101100111001111101111011111"),
                ("11111110001100111001110011100111001110011001110110100111100001000010000100001000010001011110111101111101111011010000100001000010010100101000010001001110110100111011010110101101100101100011100111011111"),
                ("11111110001100111001110011100111001110011001110110100111100001000010000100001000010001011110111101111101111011010000100001000010010100101000010001001110110100111011010110101101100101100011100111011111"),
                ("11111010001100111001110011100111001110011100110110101101101001000010000100101001010000100001000101111101101000010000100001000010011100011010110101001110110100111011010110101101100111001011000110011111"),
                ("11111110001100111001110011100111001110011100110011110100100001000010000100101000010000100001000010001011110111010000100001000010010100101001010011001110011110101001110011100111100111001110011100111111"),
                ("11111110101100111001101101011010011100111001111010010000100001001010010100101001010001101111011000011011110111101111011111011010000100101000010000100011010010011101011010100111100111001110011100111111"),
                ("11111110000110001100110011011010011100111011010110010010100101000010000100001000010000100001000010001011100001000010000110111110110100001001010010100001001100111001110011100111100111001110011100111111"),
                ("11111110000110001100110011011010011100111011010110010010100101000010000100001000010000100001000010001011100001000010000110111110110100001001010010100001001100111001110011100111100111001110011100111111"),
                ("11111010011110111101110011100110011100111011010011110100100001000010000100001000010001101111011101111011111011101111011111011010000100001000010000100011010101101011010110110011100111001110011100111111"),
                ("11111011101110111101110011100110011100111011011010010010100001000010000100001000010001101111011000011011101000010000100001000010000100001000010000100110011101101001110011100111100111001110011100111111"),
                ("11111111111111111111011001100110110101101011010011010010100001000010000100001000010001101111011110110100001000010000100001000010000100001000010000100011010100111100111001110010110010110110011100111111"),
                ("11111111111111111111111101111011001110011011010110110100100001000010000100001000010000100001000010000100001000110111101111011010000100001001010010100110011110101100011000110011110110011111111111111111"),
                ("11111111111111111111111101111011001110011011010110110100100001000010000100001000010000100001000010000100001000110111101111011010000100001001010010100110011110101100011000110011110110011111111111111111"),
                ("11111111100110001100011000110010011100111011010011100110100101001010010100101001010000100001000010001011100001101111011101000010000100011000110001001110011110100100101001100110110001110111111111111111"),
                ("11111111100110001100111101100110011100111011011010010010100101001010010100101000010000100001000110111011110111110111101101000010000100011010110101001111010101101001110011110101001101100111011110111111"),
                ("11111110011100111001110011001110110101101001101001110000100001000010000100001000010000100001000010001011110111101111011101000010000100011000110001011010011100111001110011110101001111001011000110011111"),
                ("11111100111100111001100111011010110101101001110011100110100101000010000100101000010000100001000010001011100001110111101101000010000100001001010011001110011100111001110011100111011010110011000110011111"),
                ("11111100111100111001100111011010110101101001110011100110100101000010000100101000010000100001000010001011100001110111101101000010000100001001010011001110011100111001110011100111011010110011000110011111"),
                ("11111100111011010110101101011010110101101001110110100110100101001010010100001001010000100001000010001011100001010000100001000010010100101001010010100101001100111011010110101101011010110110011100111111"),
                ("11111110011001110011100111011010011100111101010110110100100101001010010100001000010000100001000110110000110111110111101101001110000100101001010010100101001100111100111001100111100110011110011100111111"),
                ("11111111101100111001110011100110011100110100110011100111001111010110100100101000010000100001000000011011110111110111101101000010010100101001010010100101000110101100111001110011100111001110011100111111"),
                ("11111111101100111001110011100110011100111001111010100111011010011100111101001001010001011110111000011011111011010000100001000010011100001000010000100001000010011011010110100111100111001110011100111111"),
                ("11111111101100111001110011100110011100111001111010100111011010011100111101001001010001011110111000011011111011010000100001000010011100001000010000100001000010011011010110100111100111001110011100111111"),
                ("11111100111011010110101101001110110101101011010011100111011010011100111100001000010001011110111010000100001000010000100001000010011100011000110000100101000010010100101001010011100111001110011100111101"),

                -- explosion_2-2.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("10011111101111011110110011001110011100111100111110111101111111111111110111001001110001101011010110000100011000110001100001000010000100001000010000100101100111111111111111111100110011001011000110001100"),
                ("10110110011100111001100111011011001110011100101100011001111111111111111110111101011001100111001110011100111001110011100111010000111100110011100110110011110111111111111111111010110011001110011100101100"),
                ("10110110011100111001100111011011001110011100101100011001111111111111111110111101011001100111001110011100111001110011100111010000111100110011100110110011110111111111111111111010110011001110011100101100"),
                ("10110110011100111001100111011010011100111100111110011001111001100011001100111001110011011010110110011100111001101101011011010011001100111001110011100111101111101111011110011001100111001110011100111001"),
                ("10011110011100111001101101011010110101101001111001011001111011001110011100111001101101011010110110011100111001110011100111001011001001110110101101100111001110011001110011101101011010011100111001110011"),
                ("10110100111001110011100111011010110101101011010011100111100110110101101001110011100111001110011110011100111001100111001110011110101001110110101101011010110100111011010110101101011010110101101011010110"),
                ("10110100111001110011100111011010110101101011010011100111100110110101101001110011100111001110011110011100111001100111001110011110101001110110101101011010110100111011010110101101011010110101101011010110"),
                ("10110100110100101001110101001110011100111001110110101101011010110101101011010110101101001110011110011100110011101101011011010100111001110011100111011010110101101011010110100111011010110100111001110011"),
                ("10011110101001110011101101011010011100110100111010100111011010011100111101010011101101101011010100111011010110101101011010110100110100111000110001001110110101101101011010110001101010011110101101011000"),
                ("10011100111001110011110101001110011100111100001001100111101001001010010100111010010010100001000110101011010011100111001110011110100100101001010011001110011110100100101001010010100110011100111001101001"),
                ("10110101101001110011010010100101001010010100001001010010100001000010000100001000010010100001000010001101011000010010100111010010010100001000010001100001000010000100101001010011100011010110001100001000"),
                ("10011100111101011010010010100101000010000100001001010010100001000010000100001000010000100101001010000100001000010010100111000110000100001000010000100001000010000100001000010000100001001010010100101001"),
                ("10011100111101011010010010100101000010000100001001010010100001000010000100001000010000100101001010000100001000010010100111000110000100001000010000100001000010000100001000010000100001001010010100101001"),
                ("11000110100100101001010000100001001010010100001001010010100001000010000100001000010000100101001010010100101000010010100101001010000100001001010010100101001010000100001000010000100001000010000100001000"),
                ("01000010010100001000010000100101000010000100001000010010100001000010000100001000010000100101001010000100101000010000100001000010000100001000010000100001001010000100001000010000100001000010000100001000"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011011010000100001000010000100001000010000100001000010000100001000010000100011011"),
                ("10111101110100001000010000100001000010000100001000010000100011011110111101111011010001101111011010000100010111101111011100001101110000100001000011011101000010000100001000010001101101000110111101111011"),
                ("10111101110100001000010000100001000010000100001000010000100011011110111101111011010001101111011010000100010111101111011100001101110000100001000011011101000010000100001000010001101101000110111101111011"),
                ("01000000010000100001110110100001000010000100011011010000100011011110110000110111010000000100001010001011110111000010000110111101110000100001000011101101000010001011110111110111011110111000010000110111"),
                ("01000101111011110111000011011110111101111011110111101110100001000010001011110111101111011110111101111101111011101111011100001101110000100001000010100001000110111011110111101111011110111101111011111011"),
                ("01000110111011110111101110000100001000011011110111000010100001000010000100011011000011011110111101110100011011101111011100001000010000100001000010100010111000010000100001000011011100001010000100001000"),
                ("01000010001101111011110110100011011110111011111011101111101101000010000100010111000011011110111010000100001000010000100011011101110000100001000011101111011010000100001000110110000110111010000100001000"),
                ("01000010001101111011110110100011011110111011111011101111101101000010000100010111000011011110111010000100001000010000100011011101110000100001000011101111011010000100001000110110000110111010000100001000"),
                ("01000010000100001000010010100001000010000100001000010001101101000010000100011011101111101111011010000100001000010000100001000101110000110111101111011111011010000100001000010001011101000010010100101001"),
                ("01001010010100101001110000100101000010000100001000010000100001000010000100001000110110100001000010010100101001010000100001000110111011111011110110100001000010000100001000010000100001000010010100101001"),
                ("11000110000100101001010010100101000010000100001000010000100001000010000100001000010000100101001010011100001001010010100101000010000100001000010000100001000010000100001000010000100001000110101101011010"),
                ("11000010000100101001010010100101001010011100011010110000100101000010000100001000010010100001000010011101001000010000100001001010010100001000010001100001000010000100001000010000100001000010010100101001"),
                ("11000010000100101001010010100101001010011100011010110000100101000010000100001000010010100001000010011101001000010000100001001010010100001000010001100001000010000100001000010000100001000010010100101001"),
                ("01001010000100101001010010100110011100111011010011100110100101000010000100101000010000100001000100111001110011010010100101001010000100001001010011001111010010000100101001010000100001001010010100101001"),
                ("01000010000100001000010010100110011100111001111010100111001111010110101001111010010011101011010100111011010110101101011010011010000100111010110101011011010010011101011010010000100011010110101101011010"),
                ("01001010011101011010100111001110011100111001110110110101101010011100111011010110100110100101001110101001110011101101011010110100111101010011100111001111010110101001110011010010100110011110101101010011"),
                ("01001101101100111001110011011010011100111001110011010011100011001110011001110110100111101011010100111011010110101101011010011101101001111010110101011010110101101011010110010011100010011100111001110110"),
                ("01001101101100111001110011011010011100111001110011010011100011001110011001110110100111101011010100111011010110101101011010011101101001111010110101011010110101101011010110010011100010011100111001110110"),
                ("01001100111100111001100111011010011100111101011010100111100111001110011001111001100111001110011100111011010110101101011011001100111001110011100111011010110101101011010110100111101011010101101011010110"),
                ("11001110011100111001110011011010110101101001110011011001110101100011001100111001110011100111001110011100111001110011100111001011001100101100011000110011001110011011010110101101011010110101101011010110"),
                ("11001110011100111001100111011010110101101100101100011101001110110101101100111001110011100111001110011100101100110011100111001110011100111001110011111011110011000110001100011001100111001100111001111001"),
                ("11001110011100111001110011100101100011000110011101111111111111001110011100111001110011100111001110010110001110111101111011110011001100110011100111100111111111110111001110011100110011001011000110011110"),
                ("11001110011100111001110011100101100011000110011101111111111111001110011100111001110011100111001110010110001110111101111011110011001100110011100111100111111111110111001110011100110011001011000110011110"),
                ("11110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_2-3.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001111100110001100110001100001100111101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111101100110011100111001110011001110110101101011011001011000110011111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111110111001100011000110001100110011100111001110011001110110101101011010011110011100111001110011111011110111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111110111001100011000110001100110011100111001110011001110110101101011010011110011100111001110011111011110111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111100110011001110011001111001110011100111001110011001110110101101011010110101101001111001110010110001100110011111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111110111101100110011100111011010110101101011010110101101011010110100111001110011101101001111001110011100111001110011111011110111111111111111111111111111111"),
                ("11111111111111111111111111111111111111110111011110110011100110110101101011010110100111001110011100111011010110100111001111000100111011010110101101100111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111111111111111111111110111011110110011100110110101101011010110100111001110011100111011010110100111001111000100111011010110101101100111001110010110001100011001111111111111111111111111"),
                ("11111111111111111111100111100101100011000111011001110011100110110101101011010110100111011010110100111001110011110001100001000010001100010011100111011010110101101011010110011000110011111111111111111111"),
                ("11111111111111111111111100110011001110010110011001100111100110110101101011011010100111011010110110101100011000010010100101000010001100010110101101011010110101101011010110100110110011110111111111111111"),
                ("11111111111111111111111111110101100011001111001100101101001110011100111101001001110001101011010110000100101001010010100101000010000100111010110101011010110101101001110011110011110101110111101111011111"),
                ("11111111111111111111111111100111001110010110011001101101011010110101101001101001010010100101001010011100001001010010100101000010000100011000110001001110110101101001110011110010110001100111101111011111"),
                ("11111111111111111111011001100110110101101001110011101101011010110101100100101001010000100001000010000100101001010000100001000010000100011010110101001110110101101011010110110011100101100111101111011111"),
                ("11111111111111111111011001100110110101101001110011101101011010110101100100101001010000100001000010000100101001010000100001000010000100011010110101001110110101101011010110110011100101100111101111011111"),
                ("11111111111111111111110011100110110101101011010110101101011010011100110100001000010000100001000010000100001000010000100001000010000100001001010010100111010101101011010110100111100111001011000110011111"),
                ("11111111111111111111110011001110011100111011010110101101011010011100110100101000010010100001000010000100001000010000100001000010000100011000110000100111010101101011010110101101001110011110011100111111"),
                ("11111111111111111111110011001111001110011001110011100111011010011100110100101000010000100101001010000100001000010000100001000010010100101001010010100111010100111001110011110011001111001110011100111111"),
                ("11111111111111111111110011100111001110011100110011100111001111010110100100101000010010100001000010010100001000010000100001001010010100001000010000100111010110101101011010110101100111001110011100111111"),
                ("11111111111111111111110011100111001110011100110011100111001111010110100100101000010010100001000010010100001000010000100001001010010100001000010000100111010110101101011010110101100111001110011100111111"),
                ("11111111111100111001110011100111001110011100110110101101101001001010011100011000010010100001000010000100010111010000100001000010010100001000010000100110011110101101011010100111001111001110011100111111"),
                ("11111011001100111001110011100111001110011001110011110101100001001010010100101001010000100001000010001011100001101111011101000010000100001000010001001110110100111001110011101101100101100111101111011111"),
                ("11111110011100111001100111100110011100111001111010010010100101000010000100011000010000100001000010000100010111000010000110111010000100101001010011101010011100111001110011100110110001110111101111011111"),
                ("11111110011100111001101101011010110101101011011010010010100101000010000100101001010000100001000110111011110111000010000110111010000100001001010011101010011100111001110011101101100101110111101111011111"),
                ("11111110011100111001101101011010110101101011011010010010100101000010000100101001010000100001000110111011110111000010000110111010000100001001010011101010011100111001110011101101100101110111101111011111"),
                ("11111111011110111101110011001110011100111001110011100111101001001010010100001000010000100001000000011011101000110111101111011010000100101001010011100001001010011001110011100111100101100111101111011111"),
                ("11111111111111011110011001001101001010010100111010100111101001000010000100001000010000100001000000011011101000010000100001000010011100001001010010100001000010011001110011101101100101100011100111011111"),
                ("11111111111111111111011001100111010110101101011010110101101001001010010100001000010000100001000101111101101000010000100001000010000100001000010000100001000010011001110011100111100111101111101111011111"),
                ("11111111111111111111011001100110110101101011010110101101100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001110101001110011110011110101110111111111111111"),
                ("11111111111111111111011001100110110101101011010110101101100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001110101001110011110011110101110111111111111111"),
                ("11111111111111011110011001100110110101101001111010100110100101000010000100001000010000100001000010000100011011110111101101000010000100101001010010100011000010011001110011011000111011110111111111111111"),
                ("11111111101110111101110011011010110101101001111010010010100001000010000100001000010000100001000010001101100001000010000110111010000100111010110101100011010110101001110011110011100111110111101111011111"),
                ("11111111100110001100110011001110110101101011010011110000100101000010000100001000010001011110111110111011100001000010000100001010000100111000110000100111010110101001110011101101100111110111101111011111"),
                ("11111111101111011110011001100110110101101011010011010010100101001010010100001000010001101111011101110000110111101111011100001101110100010011100111001110011010011001110011101101001111001111101111011111"),
                ("11111111101111011110011001100110110101101011010011010010100101001010010100001000010001101111011101110000110111101111011100001101110100010011100111001110011010011001110011101101001111001111101111011111"),
                ("11111110011100111001110011011010110101101011010011010010100101001010010100001000010001011110111101111011101000101111011100001110110100011000110001101010011100111011010110110011100111001011000110011111"),
                ("11111111111100111001110011100110011100111101010011110100100101001010010100001000010001101111011101110000100001000010000110111010000100111000110000100111000101101011010110100111100111001110011100111111"),
                ("11111111111110111101011001111011001110011001110110110100100111000110000100001000010001101111011101111011110111101111011100001101110100010011100111001110011101101011010110100111100111001110011100111111"),
                ("11111011101111011110110011100110011100111101010011110100100101001010011100001001010001011110111101110000100001000010000110111110110100001001010011101011010101101011010110100111100111001011000110011111"),
                ("11111011101111011110110011100110011100111101010011110100100101001010011100001001010001011110111101110000100001000010000110111110110100001001010011101011010101101011010110100111100111001011000110011111"),
                ("11111011001100111001011001111011001110011001110110110100100111000110001100001001010001101111011110111011100001101111011111011010000100001000010000100110011101101011010110100111100111001011100111011111"),

                -- explosion_2-4.png
                ("11111011101100111001110011001110110101101011010011010010100001000010000100011011101110000100001101111101111011010000100001001110001100001001010011101010110100111100111001111100110011001011000110011111"),
                ("11111011001100111001110011001110110101101011011010110100100101000010001101110111000010000100001000011011110111010000100001001110000100101001010011101010011110101001110011110011100111110011100111011111"),
                ("11111110011100111001110011001110110101101011010011100111001101000010001011100001101111011110111101111011111011010000100001000010001100001001010011101010110100111100111001111100110011101111111111111111"),
                ("11111110011100111001110011001110110101101011010011100111001101000010001011100001101111011110111101111011111011010000100001000010001100001001010011101010110100111100111001111100110011101111111111111111"),
                ("11111110011100111001110011001110110101101011011000010011100001001010010100010111000010000100001000011011111011010000100001000010000100101001010011101010011110101001110011110011100111001111111111111111"),
                ("11111011001100111001110011100110110101101001110011110101100001000010001101100001101110100001000101111011110111010000100001000010000100101001010010100110011101101011010110101101100111001110011100111111"),
                ("11111111101100111001100111011010011100110100110011100111001101000010001011100001101111011110111000011011111011010000100001000010000100101001010010100110011101101011010110110010110011110111101111011111"),
                ("11111111101100111001100111011010011100110100110011100111001101000010001011100001101111011110111000011011111011010000100001000010000100101001010010100110011101101011010110110010110011110111101111011111"),
                ("11111111101111011110110011011010011100111101011010010011100001001010010100000001000010000100001101111101110111010000100001000010000100001001010011100010011101101011010110100111100101100111101111011111"),
                ("11111111101111011110110011100110011100111101011010110001101001001010010100010111000010000100001110110100001000010000100001000010000100001000010000100111010100111011010110101101100111101111101111011111"),
                ("11111111111111011110011100110010011100110100111000010000100101001010010100001000110111101111011010000100001000010000100001000010000100001001010011001111010100111011010110110010110011110111111111111111"),
                ("11111111110111001110111011100110011100111101001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110001011010110101101011010110110010110011111111111111111111"),
                ("11111111101110111101110011001110011100110100101000010000100001000010000100001000010000100001000110111011101000010000100001000010000100111010110101101011010110101101011010110010110011111111111111111111"),
                ("11111111101110111101110011001110011100110100101000010000100001000010000100001000010000100001000110111011101000010000100001000010000100111010110101101011010110101101011010110010110011111111111111111111"),
                ("11111011100110001100110011011010011100110100101000010000100111000110000100101000010000100001000101110000101000010000100001000010000100011010110101001111010010010100101001100110110011110111111111111111"),
                ("11111111100110001100110011001110011100110100101001110000100101001010010100011011110110100001000101110000101000010000100001000010000100111010110101001110011100111001110011100111100111101111011110111111"),
                ("11111111100111001110110011011010011100111001110011110100100101000010000100010111000011011110111101111101101000010000100001001010010100001001010010100111010101101011010110101101011011001110011100111111"),
                ("11111111100111001110011001001110011100111001110011110100100101001010010100010111000011011110111010000100001000010000100011000010000100001001010010100111010100111001110011110011001111001110011100111111"),
                ("11111111100111001110011001001110011100111001110011110100100101001010010100010111000011011110111010000100001000010000100011000010000100001001010010100111010100111001110011110011001111001110011100111111"),
                ("11111111100110001100110011011010011100111001110110100110100001000010000100001000101110000100001101110100001000010000100001001010010100111000110001101010011100111100111001110011100111001011000110011111"),
                ("11111110011100111001100111001111010110101101010011010010100001000010000100101000010001011110111010000100001000010010100111000110000100111010110101011010110110011100111001110011100111001111111111111111"),
                ("11111110011100111001110011101011010110101101011010010010100001000010000100101001010000100001000010000100101000010010100101000010011101010011100111001110011110011100111001110011100111111111111111111111"),
                ("11111110011100111001100111100110011100111001111010010010100101001010010100101000010000100001000010000100001001010000100001000010011001110110101101001110011100111100111001100111100111111111111111111111"),
                ("11111110011100111001100111100110011100111001111010010010100101001010010100101000010000100001000010000100001001010000100001000010011001110110101101001110011100111100111001100111100111111111111111111111"),
                ("11111110011001110011100111011010110101101011011010010011100001000010000100001000010000100001000010000100001000010010100101000010011001110110101101011010110101101001110011100111100111111111111111111111"),
                ("11111011001100111001110011001110110101101011011010010010100101000010000100001000010000100001000010000100001000010000100001000010001001110110101101011010110101101011010110110011100111111111111111111111"),
                ("11111111100110001100110011100110110101101011010110100111101001000010000100001000010000100101001010010100001000010000100001001010011011010110101101011010011100111011010110110010110011111111111111111111"),
                ("11111111100110001100011001100110011100111011010110100111100001000010000100001000010010100101001110000100101001010010100101001100111011010110101101011011001011001100111001110011111111111111111111111111"),
                ("11111111100110001100011001100110011100111011010110100111100001000010000100001000010010100101001110000100101001010010100101001100111011010110101101011011001011001100111001110011111111111111111111111111"),
                ("11111111100111001110111011100110011100111011010110101101101001001010010100001000010010100101001010011100011010110001100001001110101001110011100111011001100111100110001100111011111111111111111111111111"),
                ("11111111111111011110011001001110110101101011010110101101011011000110000100001000010011100011000110001101010110100111001111010101101011011001110011001111001011001100111001011001111011111111111111111111"),
                ("11111111111111111111011000110010110101101011010110101101001111000110000100001000110001001110011100111001110110100111001110110101101011011001110011100111001011100110001100110011001111111111111111111111"),
                ("11111111111111111111111110110001100011001100111001110011011010110101101001111000100111011010110101101001110011100111001110110101101011011001110011100111110011101111111111111111111111111111111111111111"),
                ("11111111111111111111111110110001100011001100111001110011011010110101101001111000100111011010110101101001110011100111001110110101101011011001110011100111110011101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111110111101100111001110011100110011100111011010011100111011010110101101011010110101101011010110101101001111001110011111011110111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111100101100011001100110011100111011010110101101011010110100111100111001110011100111001100111100101100011001111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111110111101100111001110011100110011101101011010110100111100111001110011100101100011000110001110011101111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111101100011000110011001101101011010110100111100111001110011100101100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111101100011000110011001101101011010110100111100111001110011100101100111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111001100110000110001100011001111011001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_2-5.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("01100011101111111111111111100111110111101111011110111111111111111111111111111101110011100111001011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11001111101110111101110011100111110111100110011101111101111111111111111111011101110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11001111101110111101110011100111110111100110011101111101111111111111111111011101110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("01100110010110001100110011100101100011001100111001011000110001100011000110011001101101001110011110011100111001110011100111001110010110011111111111111111110100111111111111111111111111111111111111111111"),
                ("11110110011111011110110011011011001110011001110110110011100111001110011001110011101101100111001110011100111001100111001110011110011100111001110011110101100110011111111111111111111111111111111111111111"),
                ("11001100111100111001100111011010110101101011010110101101011011010110100100110011101101001110011110011100111001110011100110011101101011011001110010110011001011001111111111111111111111111111111111111111"),
                ("11001100111100111001100111011010110101101011010110101101011011010110100100110011101101001110011110011100111001110011100110011101101011011001110010110011001011001111111111111111111111111111111111111111"),
                ("10011110101001110011110101011010110101101011010011100111011011010110100100110011101101001110011100111100111001100111001110110101101001101100011001111001100011100111001110111111111111111111111111111111"),
                ("10110100111011010110100111001110011100111001111010110101011011010110101101010011110101101011010100111011010011100111001110110101101001111001110010110011001110011111011110111101111111111111111111111111"),
                ("11010110101101011010110100100101001010011100001001100111011011010110101001110011010010100101001110101011010011100111001110110101101011010110101101011010011110011100111001111101111011111111111111111111"),
                ("01001010010100101001010010100101001010010100101000010011100011010110101101011010010010100101001110001101010011101101011010110101101011010110101101001111001110011100111001110010110001110111111111111111"),
                ("11000010011100011000010010100101001010010100001000010000100001001010010100001001010000100001000010010100111010100111001110011100111011010110101101001110110101101011010110100111100101100111111111111111"),
                ("11000010011100011000010010100101001010010100001000010000100001001010010100001001010000100001000010010100111010100111001110011100111011010110101101001110110101101011010110100111100101100111111111111111"),
                ("11000110000100001000010000100001000010000100001000010000100001000010000100001000010010100001000010011100001001010010100101001010000100110011100111101010110101101011010110101101001101100111111111111111"),
                ("01001010010100001000010000100001000010000100001000010000100001000010000100001000010011100011000010011100001000010000100001000010000100101001010010100111010101101011010110101101100101100011000110011111"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010000100001001010000100001001010011100010011100111001110011101101100111001110011100111001"),
                ("11011101111101111011110111011111011110111011101000010000100001000010000100001000010000100001000010000100001000010010100101000010000100001001010011101010110101101001110011101101100111001110011100111001"),
                ("11011101111101111011110111011111011110111011101000010000100001000010000100001000010000100001000010000100001000010010100101000010000100001001010011101010110101101001110011101101100111001110011100111001"),
                ("11011101111011110111101111011110111101111101101000010000100010111101110000100001110110100001000010000100001001010000100001000010000100001001010011100011010100111001110011101101100111001110011100111110"),
                ("10111000011011110111000011011100001000011011111011010000100011011110111011110111101110100001000101110100001000010000100001000010000100111000110000100111000100111011010110101101001110011100111001101100"),
                ("00001000011011110111000010100010111101110000100001110110100001000010000100001000101111011110111000011011101000010000100001000010000100101001010010100111000100111011010110101101011010110101101011001100"),
                ("10111000011011110111000011011110111101110000100001110110100001000010000100011011000010000100001101110100001000010000100001000010000100001001010010100101001110001001110011100111011010110101101011011000"),
                ("10111000011011110111000011011110111101110000100001110110100001000010000100011011000010000100001101110100001000010000100001000010000100001001010010100101001110001001110011100111011010110101101011011000"),
                ("11011101110000100001101110000100001000010000110111010000100001000010000100011011101111011110111010000100001001010000100001000010000100001000010000100001000010001100011000100111011010011110011100101100"),
                ("01000110111011110111010001101110111101110100001000010000100001000010000100101000010000100001000010000100101001010010100101000010000100001000010000100001000010001001110011101101011011001011000110011110"),
                ("01000010000100001000010010100001000010000100101001010010100001000010001100001001010000100101001010000100001000010010100101000010000100001000010000100111000110001011010110100111001111001011000110011111"),
                ("01000010011001110011110001100010011100111100011010010010100001000010000100101001010010100101001010000100001000010010100111000010011101011000110001101010110100111011010110110011100111001111111111111111"),
                ("01000010011001110011110001100010011100111100011010010010100001000010000100101001010010100101001010000100001000010010100111000010011101011000110001101010110100111011010110110011100111001111111111111111"),
                ("01001110101001110011010011101010011100110100111000010000100001000010000100011000110101101011010100110100101001010010100101001010011001110011100111011010110101101100111001110010110011110111111111111111"),
                ("10011110101001110011110001001110011100111101011010110000100101000010000100001001100111001110011101101001111010110101101011010110101011010110101101011010110101101100111001110010110011110111111111111111"),
                ("10110101101011010110101101001101001010011101011010010011101001001010010100101001100111001110011100111101011010100111001110110101101011010110101101011010110101101100111001110011100111111111111111111111"),
                ("10110101101011010110101101011010011100111001110011100111001110011100111001110011100111001110011100111101011010100111001110110101101011010011100111001110110101100110001100111101111111111111111111111111"),
                ("10110101101011010110101101011010011100111001110011100111001110011100111001110011100111001110011100111101011010100111001110110101101011010011100111001110110101100110001100111101111111111111111111111111"),
                ("10011100111001110011100111100110110101101011011001011001100110011100111011010011101101001110011101101001111010110011100110110100111100111001110011100110011011000110001100111111111111111111111111111111"),
                ("11001110011100111001110011100110011100111100111001011101110111001110011100111001110010110001100110011001111001100111001110011110011100101100011001110101100011001111111111111111111111111111111111111111"),
                ("11001110011100111001110011100111001110011111011110111100111011101111010110001100011100111001110011001100111001110011100110011110010110001100011000111011110111111111111111111111111111111111111111111111"),
                ("01110011001100111001110010110011110111101111011110111111111111110111100111011110111101111011110111101100111001110011100111001011001111011110111101111011111111111111111111111111111111111111111111111111"),
                ("01110011001100111001110010110011110111101111011110111111111111110111100111011110111101111011110111101100111001110011100111001011001111011110111101111011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_2-6.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111101111011110111100110011001110011100111001110011111011110111101111011110011101111011111111111111111110111101111011110011001100111001011000110001110"),
                ("11111111111111111111111111111111111111111111111110011100110001100011001100110011110011100111001110010110001110011100111001100011001110101110011101111011110111101100111001110011100111001110011100111001"),
                ("11111111111111111111111111111111111111111111111110011100110001100011001100110011110011100111001110010110001110011100111001100011001110101110011101111011110111101100111001110011100111001110011100111001"),
                ("11111111111111111111111111111111111111110110001100111010110011001110011100110011100111100111001100111100101100110011100111001110011100111101111010111011001110011001110011110011100111001110011100111001"),
                ("11111111111111111111111111111101100011000110010011110011100111001110011001110110110011101011010100111011010011101101011010011101101001111001110010110011001101101011010110110011001110011100111001110011"),
                ("11111111111111111111111111111001100011001011010110100111001110110101101011010110100111101011010110101001110011100111001110011100111001110011100111001110011100111001110011101101011010110101101011010110"),
                ("11111111111111111111111111111001100011001011010110100111001110110101101011010110100111101011010110101001110011100111001110011100111001110011100111001110011100111001110011101101011010110101101011010110"),
                ("11111111111111111111110011100111001110011011010110101101011010110101101011010110100111101011010110101001110011100111001101001010010100111010110100100111010110100100101001100111011010110101101011010110"),
                ("11111111111111011110011001100111001110011011010110101101011010110101101101011010110101101011010100111011010011100111001101001010000100001001010011100011010110101001110011100111100010011110101101010011"),
                ("11111111111111011110011001100111001110011011010110101101001110011100110100101001010010100101001010011001111010110101101011000010000100001000010000100011000010011001110011110100100110011110101101001001"),
                ("11111111111100111001110011100110110101101001110110110101100011010110100100111000010010100001000010000100001001010010100101001010010100001000010000100111010110001001110011110001100010011010010100101000"),
                ("11111011001100111001100111001110110101101100011000010010100001000010000100001000010010100001000010000100001001010000100001001110000100001000010000100101001010010100001000010000100101000010000100001000"),
                ("11111011001100111001100111001110110101101100011000010010100001000010000100001000010010100001000010000100001001010000100001001110000100001000010000100101001010010100001000010000100101000010000100001000"),
                ("11110011001100111001101101011010011100110100001000010000100001000010000100001000010010100101001010010100001000010000100001000010010100001000010000100001000010001011110111110110100010111110111101101000"),
                ("01100110011001110011101101001111000110000100001000010000100001000010000100001000010000100101001010000100010111101111011111011010000100001000010000100010111000010000100001000011011100001101111011111011"),
                ("11000101101011010110101101001110011100111100001001010010100101000010000100001000010000100001000010001011100001000010000111011010000100001000010001101100001000011011110111101110000110111000010000110111"),
                ("01100101101011010110101101011010110101101001111000010010100101001010010100001000010000100001000101110000110111101111011101000010000100001000010001101100001000011011110111010000000110111000010000100001"),
                ("01100101101011010110101101011010110101101001111000010010100101001010010100001000010000100001000101110000110111101111011101000010000100001000010001101100001000011011110111010000000110111000010000100001"),
                ("01100100111001110011100111011010110101101001111000010011100001001010010100001000010000100001000010001011101000101111011110111101111101101000010000100011011101110000100001101110000110111000010000110111"),
                ("11110110011100111001110011011010011100111001111010110000100101000010000100001000010000100101001010000100001000110111101100001000011011101000010000100001000110111011110111101111011110111101111011111011"),
                ("11001110011100111001110011011010011100111011010110110100100101000010000100001000010010100001000010000100001000010000100001000010000100001000010000100001000101111101111011101111101111011101111011111011"),
                ("11001110011100111001110011011010011100111001110011110000100101000010000100001001010000100101001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("11001110011100111001110011011010011100111001110011110000100101000010000100001001010000100101001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("11111011000110001100110011011010110101101011011010010010100101001010010100001000010000100001000110000100111000010010100101000010000100001000010000100001000010000100001000010000100001000010010100101001"),
                ("11111111110110001100100111011010110101101011010110110101001101001010010100001001010010100101001110000100101000010010100101000010000100001000010000100001000010000100001000010000100001000110001100011000"),
                ("11111111110110001100110011001110110101101011010110100111011010110101101001110011100111101011010010010100101000010000100001001010000100101000010000100001000010000100101001010010100111000010010100111000"),
                ("11111111110111001110011001100111001110011100111001100111011010110101101011010110101101001110011110101100001001010010100111010110101101011000110000100101000010010100101001010010100101001010010100101001"),
                ("11111111110111001110011001100111001110011100111001100111011010110101101011010110101101001110011110101100001001010010100111010110101101011000110000100101000010010100101001010010100101001010010100101001"),
                ("11111111111111111111111101111011001110011100110011101101011010110101101011010110100111001110011101101101001001010010100110011100111101010110101101001101001110000100101001010011101011010110101101011010"),
                ("11111111111111111111111111111011110111101100111001011001100110011100111011010110100111001110011101101001111010110101101010011110101101010110101101101011010100111001110011100111001110110100111001110110"),
                ("11111111111111111111111111111101110011100111001100111100110010011100111011010110100111100111001110011001110011101101011010011010011101010110101101001110011101101011010110101101101010011110101101010011"),
                ("11111111111111111111111111111111111111110110011001011001100110110101101011010011110011100111001110011100110011101101011010011010011101010110101101011010110101101011010110101101001111001100111001111001"),
                ("11111111111111111111111111111111111111110110011001011001100110110101101011010011110011100111001110011100110011101101011010011010011101010110101101011010110101101011010110101101001111001100111001111001"),
                ("11111111111111111111111111111111111111111100101100111011100111001110011100110011100111100111001110011100111001101101011010011100111100111001110011100110110100111100111001101101100111110110011100111110"),
                ("11111111111111111111111111111111111111111001111110111111111101100011001100111001110011100111001110011100110011101101011011001011000110001100011000110011001110010110001100110011100101100110011100101100"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111101111101111111111111111111011101011001111011110110011100111101111101111011001"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001110011100111101111111111111111111111111111110111101111011110110011111111111011100111001100"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011001110011100111101111111111111111111111111111110111101111011110110011111111111011100111001100"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_3-0.png
                ("11111111111111011110111100110001100011001011001001010000100001000010001101100001000010000100001000010000110111101111011111011010000100101001010010100111010101101001110011110010110001110111111111111111"),
                ("11111100111100111001110011100111001110011001101001010000100001000010000100011011101111011110111000010000100001000010000100001010000100001000010000100001001110101101011010100111001101100100111001110011"),
                ("10110100111100111001110011001110011100110100101001010000100001000010000100001000010000100001000000010000100001101111011101000110110100011000110000100001000010011101011010110101101010110101101011011001"),
                ("10110100111100111001110011001110011100110100101001010000100001000010000100001000010000100001000000010000100001101111011101000110110100011000110000100001000010011101011010110101101010110101101011011001"),
                ("10110101101100111001110011001110011100110100101000010000100001000010000100001000010001011110111000011011111011010000100001000101110000101001010010100101001110101101011010010010100110011100111001110011"),
                ("10011101101011010110100111101001001010010100101000010000100001000010000100011011101111011110111000011011110111010000100001000101110000110111101110100011000110001100011000010010100101001010010100111010"),
                ("10011101101001110011110100100101001010010100101001010000100001000010001011100001000010000100001000010000100001101111011110111101111011101000010000100011000010010100101001010010100001000010000100001001"),
                ("10011101101001110011110100100101001010010100101001010000100001000010001011100001000010000100001000010000100001101111011110111101111011101000010000100011000010010100101001010010100001000010000100001001"),
                ("10110100111001110011110100100101001010010100001001010010100011011110110000100001000010000100001000010000100001000010000100001000010100001000010000100001001110000100101001010000100001001010010100101001"),
                ("11010110100100101001010010100101000010000100001000010001101100001000010000100001000010000100001000010000100001000010000100001000010100011011110110100001001110000100101001010010100101001110001100011000"),
                ("01001110100100101001010010100101000010000100001000110111011111011110111011110111000010000100001000010000100001000010000100001101111011110111101110100001001110001100011000010010100101001010000100000011"),
                ("10011110100100001000010000100111011110110100001000010001011111011110110100010111000010000100001000010000100001000010000100001101110000100001000010100001001110000100001000010000100001000010000100001110"),
                ("01001010000100001000010000100001000010000100001000010001011111011110110100010111000010000100001000010000100001000010000110111101111011100001000010100001000010010100001000010001101110111110101101011001"),
                ("01001010000100001000010000100001000010000100001000010001011111011110110100010111000010000100001000010000100001000010000110111101111011100001000010100001000010010100001000010001101110111110101101011001"),
                ("01001010011101111011101110100011011110111101110111110110100011011110110000100001000010000100001000010000100001101111011101000010000000100001000011101110111101110100001000010000000100001101111011111000"),
                ("01001010001101111011010000100011011110111011100001000011011110111101110000100001000010000100001000010000100001000010000101000010000000100001000011101110111000011011110111101111011100001101111011100001"),
                ("01000110111011110111010000100010111101110000110111000010000100001000010000100001000010000100001000010000100001101111011101000110111101100001000011011111011000010000100001110110100011011101111011100001"),
                ("01000101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000101000000010000100001101111101101000110111101100001"),
                ("01000101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000101000000010000100001101111101101000110111101100001"),
                ("00001000011011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111011000010000100001000011011101000110111101100011"),
                ("10111000011011110111101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110111101111011101100"),
                ("01000110110000100001101111011100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011"),
                ("01000010001101111011101110000100001000010000110111101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001101110000100001000010000100001"),
                ("01000010001101111011101110000100001000010000110111101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001101110000100001000010000100001"),
                ("01000010001011110111101111011111011110111011110111010000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001101111101111011110111101110111000010000100001"),
                ("11011010000100001000010000100010111101110000110111101110000100001000010000100001000010000100001000010000100001000010000100001000011011110111101111101110111101111011110111010000100001000110111101110111"),
                ("01000010000100001000010000100010111101111011101000101111011100001000010000100001110111011110111000010000100001000010000100001000010100001000010000100010111101111101111011010000100001000010000100001000"),
                ("01000010000100001000010000100001000010001010101001110111011110111101111011111011000010000100001000010000100001000010000100001101111101110111101110100010111101110100001000010000100001000010000100001000"),
                ("01000010000100001000010000100001000010001010101001110111011110111101111011111011000010000100001000010000100001000010000100001101111101110111101110100010111101110100001000010000100001000010000100001000"),
                ("01001010000100001000010010100001000010000100001001010000100001000010000100010111000010000100001000010000100001000010000110111010001011110111101110100001000010000100001000010000100001000010010100111110"),
                ("11000110000100101001010000100101001010010100101000010000100001000010001101110111000010000100001101111101101000101111011100001000010000111011110110100001000010000100001000010000100101001010000100001001"),
                ("01001010010100101001010011101010011100111100001001010000100010111101111011110111101111011110111101111101101000101111011100001000010000110111101110100001000010000100001000010010100111000010000100001000"),
                ("01001010010100101001010011001110011100111100001001010000100010111101110100010111000011101111011010000100001000101111011100001101111011101000010000100101001010000100001000010010100101001100111001111010"),
                ("01001010010100101001010011001110011100111100001001010000100010111101110100010111000011101111011010000100001000101111011100001101111011101000010000100101001010000100001000010010100101001100111001111010"),
                ("11000110001100011000110101011010011100110100101000010000100001000010000100010111000010000100001101111011110111101111011100001101110100001000010001101011000010010100101001010011100010011100111001110011"),
                ("11001011001001110011110100100111010110101101001000010000100001000010000100010111000010000100001000010000110111101111011100001101110100001000010000100101000010011101011010110001001110011110011100111001"),
                ("11110111101001110011010010100101001010010100101001010010100101000010001101100001000010000100001000010000110111000010000110111101110100001000010000100001000010010100101001010011101011001110011100111101"),
                ("11111111011100111001100110100101001010010100001001010010100010111101110000100001000010000100001000010000100001000010000110111101110100001000010000100001001110000100101001110101001111001110011100111111"),
                ("11111111011100111001100110100101001010010100001001010010100010111101110000100001000010000100001000010000100001000010000110111101110100001000010000100001001110000100101001110101001111001110011100111111"),
                ("11111111111100111001100110100001000010000100001001010001011100001000010000100001000010000100001000010000100001000010000100001000011101101000010000100001001010011001110011110011100111001111111111111111"),

                -- explosion_3-1.png
                ("10110100111001110011101101011010110101101011010110101101001101001010010100001000010000100001000010000100001000010000100001000010010100111010110100100001000010000100101001100111001111001011000110001100"),
                ("01100110011100111001100111001110110101101001110011100111101001001010010100011011101110000100001110110100001000110111101111011010000100001000010000100001000010000100001000010010100110011110011100111001"),
                ("11101111100110001100100111011010011100110100101000010000100001000010001101100001000010000100001110110100010111000010000110111010000100001000010000100101000010010100101001010011101011001110011100111111"),
                ("11101111100110001100100111011010011100110100101000010000100001000010001101100001000010000100001110110100010111000010000110111010000100001000010000100101000010010100101001010011101011001110011100111111"),
                ("11111111110110001100110011100110011100110100101000010000100001000010001010110111000011011110111101111011100001000010000110111110110100101001010010100101000110001101011010110101001111001111111111111111"),
                ("11111111111110111101110011100111010110100100101001010000100001000010000100001000101111101111011000010000100001000010000100001101110100001000010000100101000110001001110011101101001111001111111111111111"),
                ("11111111111100111001101101100111010110100100001001010010100101001010010100001000101110000100001000010000110111000010000100001000011101101000010000100101001110001011010110110011100111001011000110011111"),
                ("11111111111100111001101101100111010110100100001001010010100101001010010100001000101110000100001000010000110111000010000100001000011101101000010000100101001110001011010110110011100111001011000110011111"),
                ("11111111110110001100101101011010011100110100001001010000100101001010010100111011101110000100001110111011110111000010000100001000011011101000010000100001001110001001110011101101001111001111101111001110"),
                ("11111111111001110011101101011010011100110100111000010010100101000010000100001000000011011110111110110000100001000010000110111101110100001000010000100001001010011001110011101101011011001011000110001100"),
                ("11111111111011010110101101011010011100110100101001110000100101000010000100001000110110000100001000011011100001000010000110111010000100001000010000100001000110101011010110101101011010110100111001111001"),
                ("01100101101001110011110101001111010110101100001001010010100101000010000100011011101110000100001000011011111011000010000110111010001101101000010000100001000010011001110011100111001111001110011100111001"),
                ("11001100111001110011110100100101001010010100101000010000100001000010000100010111000010000100001000011101101000101111011100001000011011101000010000100001000010000100101001110101100111001110011100111111"),
                ("11001100111001110011110100100101001010010100101000010000100001000010000100010111000010000100001000011101101000101111011100001000011011101000010000100001000010000100101001110101100111001110011100111111"),
                ("11001110011011010110100110100101001010010100001000010000100001000010000100010111000010000100001000010000100001000010000110111010000100001000010000100001000010011101011010101101011010110111111111111111"),
                ("11010110011011010110110100100111000110000100001000010010100001000010001101100001000010000100001000011011100001101111011100001110110100001000010000100001001010011101011010101101011010110111111111111111"),
                ("11001110011011010110100111101010011100111100001001010010100001000010001101100001000010000100001000011011100001010000100011011110110100001000010000100001001110001001110011101101011010110111111111111111"),
                ("10110110011100111001101101011010110101101101001000010010100001000010000100011011000011011110111101111011110111101111011101000010000100001000010000100101001010011101011010110101001110110111111111111111"),
                ("10110110011100111001101101011010110101101101001000010010100001000010000100011011000011011110111101111011110111101111011101000010000100001000010000100101001010011101011010110101001110110111111111111111"),
                ("01100100111100111001101101011010011100111100001001010010100111011110111011111011101110100001000010000100011011101111011111011010000100001000010000100101001010011101011010110101001110011110011100111101"),
                ("11001100111011010110100111011010110101101101001000010000100001000010001101101000010000100001000010001101110111110111101101000010000100001000010000100001000010001101011010100111011011001011000110001100"),
                ("11001110011100111001110011001110110101101101001000010000100001000010000100001000010001011110111110111011110111101111011101000010010100001000010000100001000010011001110011100111100101100011000110011001"),
                ("11010011001100111001110011011010011100111101001001010000100001000010000100011011101110000100001000010000111011000010000101000010010100101000010000100001000010011001110011100111001111110011000110011111"),
                ("11010011001100111001110011011010011100111101001001010000100001000010000100011011101110000100001000010000111011000010000101000010010100101000010000100001000010011001110011100111001111110011000110011111"),
                ("11111111111100111001110011011010110101100100101000010000100001000010001101100001000010000100001000011101111011000010000111011010000100001001010010100101001010001101011010100111001110011111111111111111"),
                ("11111111111100111001100111001110011100110100001000010000100001000010000100001000101111011110111110111101110111000010000110111010000100001000010000100111000110101100011000100111001111001111111111111111"),
                ("11111111111101011010110000100101000010000100001001010000100001000010000100001000110111101111011101110000100001000010000110111010000100101001010011100001001010011100011000100111001111001011000110011111"),
                ("11111111110100101001010010100101000010000100001000010000100001000010001011110111101111011110111000010000100001101111011111011010000100101001010011100011000010011001110011110011100111001110011100111001"),
                ("11111111110100101001010010100101000010000100001000010000100001000010001011110111101111011110111000010000100001101111011111011010000100101001010011100011000010011001110011110011100111001110011100111001"),
                ("11111111111001110011100111001111010110100100001000010000100001000010001101100001000011011110111000011011110111110111101111011010000100001000010000100101001110101001110011101101001111001110011100111001"),
                ("11111111111011010110101101011010011100111100001001010000100001000010001101100001000010000100001000011101101000101111011110111010000100001000010000100001000010011011010110101101001111001110011100101100"),
                ("00011011001011010110101101011010110101101001101001010000100001000010001011100001000010000100001000010000100001110111101100001110110100001000010000100001000010001001110011101101011001100111101111011110"),
                ("11010111011011010110101101001110110101101101001001010000100001000010000100010111000010000100001000010000100001110111101100001110110100001000010000100001000010011011010110100111011011110111101111001100"),
                ("11010111011011010110101101001110110101101101001001010000100001000010000100010111000010000100001000010000100001110111101100001110110100001000010000100001000010011011010110100111011011110111101111001100"),
                ("11001110011011010110100111001110011100111100001000010001101110111101111011100001000010000100001000010000100001101111011110111010000100001000010000100001000010001001110011100111001101100111111111111111"),
                ("11001110011001110011101101011011000110000100101000010001101100001000010000100001110111011110111000010000100001000010000100001101110100001000010000100001000010001100011000100111100111101111111111111111"),
                ("11110111011100111001101101001101001010010100001001010000100011011110110000100001101110000100001110110000100001000010000100001101111011101000010000100001001010011001110011100110110001110111111111111111"),
                ("11111011100110001100110011001101001010011101001001010000100001000010001011100001101111011110111110110100000001101111011101000010000100001000010000100001001110001101011010100111100111001111111111111111"),
                ("11111011100110001100110011001101001010011101001001010000100001000010001011100001101111011110111110110100000001101111011101000010000100001000010000100001001110001101011010100111100111001111111111111111"),
                ("11111111110110001100111010110011010110101001101001010000100001000010001011111011010001101111011110110100010111101111011101000010000100001000010000100001001110000100101001110001001110110111111111111111"),

                -- explosion_3-2.png
                ("11111111111111011110110011100111010110100001111111111111111111111111111111111111110101100111001110010110010110110011100111010110011100101100011001111111111111111111111111111111111111101011000110010110"),
                ("11111011101110111101110011100111101111010110011111111111111111111111111111111111011001100111001100111001111001110011100111001110011001110110101101111111111111111111111111111111111111110110011100110011"),
                ("01100011001100111001100111011010110101101011010110100110100111010110101100111001110011100111001101101100111001101101011010110101101001110011100111011010011011001100111001111010110001100110011100110011"),
                ("01100011001100111001100111011010110101101011010110100110100111010110101100111001110011100111001101101100111001101101011010110101101001110011100111011010011011001100111001111010110001100110011100110011"),
                ("11101110011011010110101101001110110101101011010110100110100111000110001001111001110011100111001100111011010110100111001111010100111101011010110101011010110101101011010110110011100110011100111001110110"),
                ("01100100111001110011101101001110011100111011010110100110100101001010011001110110101101001110011101101011010110110101101001001010010100110011100111011010110101101100111001110011100110110100111001110110"),
                ("11010010010100101001110001001110110101101011010011110100100001000010001001110110100111011010110101101001110110100111001111000010010100111010110101001110011100111101011010110101001110011101101011010110"),
                ("11010010010100101001110001001110110101101011010011110100100001000010001001110110100111011010110101101001110110100111001111000010010100111010110101001110011100111101011010110101001110011101101011010110"),
                ("10011110100100001000010011100011010110101001111000010000100001000010000100001001110101101011010110101100011010110001100001000010000100111000110000100101001010000100001000010010100101001100111001110110"),
                ("01001010010100101001010000100001001010010100101001010000100001001010010100001000010010100001000010000100101000010010100101000010000100001001010010100111000010010100101001010010100001000100111001110110"),
                ("01000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010000100001001010011100001001010000100101001010000100001000100111001110110"),
                ("01000010000100001000110111101101000010000100001000010000100001000010000100001000010000100001000010000100101000010000100001000010000100001001010010100101001010010100101001010000100001000110101101010011"),
                ("01000010001101111011000011011101000010000100001000010000100001000010000100001000010000100001000010001101101000010000100001000010000100001000010000100001000010010100101001010000100001000010010100101001"),
                ("01000010001101111011000011011101000010000100001000010000100001000010000100001000010000100001000010001101101000010000100001000010000100001000010000100001000010010100101001010000100001000010010100101001"),
                ("10111101110000100001000011011101000010001011111011110111011101000010000100011011010000100001000110111011101000110111101111011010000100001000010000100001000010010100001000010001010111011010000100001000"),
                ("11011000010000100001000010000110111101110000100001000011011101000010000100000001110110100001000010001101111011000010000100001101111011111011110110100001000110110100001000010001011100001110111101101000"),
                ("01000101111011110111110110000100001000010000100001000011011111011110111011100001101110100001000010001011100001000010000100001000010000110111101111101100001101111011110111101110000100001101111011101000"),
                ("11011101110000100001101110000100001000010000100001101111011111011110111011100001000011011110111010000100010111000010000100001000010000100001000010000110111000010000100001110111011100001000010000101000"),
                ("11011101110000100001101110000100001000010000100001101111011111011110111011100001000011011110111010000100010111000010000100001000010000100001000010000110111000010000100001110111011100001000010000101000"),
                ("11011110111101111011000010000100001000010000100001000010000110111101111101100001000011101111011010000100010111000010000100001000010000100001000010000111011110110000100001000011011111011110111101101000"),
                ("01000010000000100001000010000100001000010000111011101110000100001000011101111011000011011110111110110100010111101111011110111000011101110111101111011100001101110000100001000011011101000010000100001000"),
                ("10111000010000100001000010000100001000010000101000101110000100001000011011111011110111011110111101111101110111000010000100001000010100011011110110000100001101111011110111000010000110111010000100001000"),
                ("10111101110000100001000011011111011110111101110111110111011100001000010000100001000011011110111110111011110111010000100010111000011011100001000010000100001000010000100001000010000100001110111101101000"),
                ("10111101110000100001000011011111011110111101110111110111011100001000010000100001000011011110111110111011110111010000100010111000011011100001000010000100001000010000100001000010000100001110111101101000"),
                ("01000010000000100001000011011100001000010000110111110111101110111101111011111011010000100001000010001101101000110111101100001101110000110111101111011110111000010000100001000011011110111110111101101000"),
                ("01000010001011110111101110100011011110111101101000010000100001000010000100001000010010100101001010000100001000110111101111011010000000101000010000100010111000010000100001101111101101000010000100001001"),
                ("01000010001011110111010000100001000010000100001000010000100101001010010100001000010010100001000010000100001000010000100001000010001011111011110110100001000101111101111011010000100101000010000100001001"),
                ("01000010000100001000010000100001000010000100001000010000100101001010010100001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101000010000100011010"),
                ("01000010000100001000010000100001000010000100001000010000100101001010010100001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101000010000100011010"),
                ("01000010000100001000010000100001000010000100001000010011100011000110000100101001010000100001000010000100101001010000100001000010000100001000010000100001000010000100101001010010100101001010000100001000"),
                ("01001010010100101001010000100001000010000100001000010011100001001010011100001001010000100001000010000100101001010010100101001010000100001000010000100001001010010100101001010000100001000010000100001000"),
                ("11000110000100101001010000100001001010010100001001110100100101001010011101001000010010100101001010000100101001110001100001001010010100001001010011101001001110001100011000110001100001001010000100001000"),
                ("01001110101001110011110001001110110101101001110110100111001111000110001100011010100111001110011110101101011010100111001111010110100100110011100111011010011100111011010110100111101001001010000100001001"),
                ("01001110101001110011110001001110110101101001110110100111001111000110001100011010100111001110011110101101011010100111001111010110100100110011100111011010011100111011010110100111101001001010000100001001"),
                ("11000100111001110011100111001110011100111011010110101101100110011100111001110011100111001110011100111101011010101101011010110101101101010011100111011010110101101100111001101101101001001010010100110011"),
                ("10011110010110001100110011001110110101101011010011100111100110011100111001110011100111100111001101101001110011101101011010110101101100110011100111011010110100111100111001100111001111010010010100110011"),
                ("10110110010111001110111010110011110111100110011001110011100111001110011100110011111100110001100110011001110110101101011010110101101100111001110011011011001110011100111001110011100111001100111001111001"),
                ("11111111111111111111111111111111110111101111011001110011100101100011001111111111011000110001100011001100111111111111111111111111111100111001110011001101100111100110001100111111111111001110011100101100"),
                ("11111111111111111111111111111111110111101111011001110011100101100011001111111111011000110001100011001100111111111111111111111111111100111001110011001101100111100110001100111111111111001110011100101100"),
                ("11111111111111111111111111111101100011001111001100110011100111111111111111111111111111100111001011001110111111111111111111111111111111111001110011100101100011101111111111111111111111111110011100101100"),

                -- explosion_3-3.png
                ("11001111111111111111111111111111111111111111111111111111110111001110011100111001110011001110011100111001111001100111001101001010010100111010110101111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111100111001110011001110011100111011010110101101011011001100111001110011100111101001100011001111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111011010110110011100110110101101011010110101101011010110101101011010110100111001111001110011100101100011000110011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111011010110110011100110110101101011010110101101011010110101101011010110100111001111001110011100101100011000110011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111110110101101011010110101101001110011100111011010110101101011010110101101011010110100111001110011100111011010011100111001110011111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111011010110101101011010011110100100111010110101011010110100111001110011101101001110110101101011010011101101101011010110101011001100111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111001111010110101001110011010010100111010110101001110110100111001110011101101101011010110101101010011101101001111000110001001110110011000110001100111111111111111111111111111111"),
                ("11111111111111111111111111001111010110101001110011010010100111010110101001110110100111001110011101101101011010110101101010011101101001111000110001001110110011000110001100111111111111111111111111111111"),
                ("11111111111111111111111111101001001010011101011010010011100001001010011100001001100111011010110100111100001001110001100010110101101101001001010011101010110110011100111001011101111111111111111111111111"),
                ("11111111111111111111101101101001001010011100001000010000100001000010000100101001110001001110011110000100101001010010100110011101101101001001010011100010011100110110001100111101011011111111111111111111"),
                ("11111111111100111001101101101001001010011100001001010000100001000010000100001001110001101011010010010100101000010000100001000010010100101001010011100001001110101100111001101101011001100111111111111111"),
                ("11111111111001110011100111100001001010010100101001010000100101001010010100001000010010100101001010010100001000010000100001000010000100001001010010100101001100111011010110101101011011001111111111111111"),
                ("11111111110110001100110011101001001010010100101000010000100101001010010100101000010000100001000010010100001000010000100001000010000100101001010010100010011101101001110011110010110001100111111111111111"),
                ("11111111110110001100110011101001001010010100101000010000100101001010010100101000010000100001000010010100001000010000100001000010000100101001010010100010011101101001110011110010110001100111111111111111"),
                ("11111111111111011110110011001111010110100100101001010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100111010101101011010110110011100101100111111111111111"),
                ("11111111111110111101110011011011010110100100101000010000100101001010010100001000010000100001000010000100001000110111101101000010000100001000010000100111010101101011010110101101011011001111111111111111"),
                ("11111111101111011110100111011011010110100100101001010000100001000010000100001000010000100001000010000100011011110111101101000010000100001000010000100011010101101011010110101101011011001111011110111111"),
                ("11110011001110111101101101011010011100111100001001010010100001000010000100010111101111101111011010000100010111110111101101000010000100001000010000100001000110001101011010110101001110011011000110001100"),
                ("11110011001110111101101101011010011100111100001001010010100001000010000100010111101111101111011010000100010111110111101101000010000100001000010000100001000110001101011010110101001110011011000110001100"),
                ("11110110011100111001011001011010110101101011011010010010100101000010000100010111000011011110111000010000110111101111011101000010000100001000010000100001000010000100101001010011101011010110011100111001"),
                ("11001110011100111001100111001110110101101011011010010000100001000010000100010111000011011110111101111011100001101111011101000010000100001000010000100001000010000100101001010011101010011110011100111001"),
                ("11001011001111011110111101100111001110011011011010010000100001000010001101100001101110000100001101111101111011000010000111011010000100001000010000100001000010000100101001110001001110011110011100111001"),
                ("11111011000111001110111100110011001110011011010011010000100011011110110000100001101111011110111101110000101000101111011110111010000100001001010010100001000010011101011010100110110001100110011100111111"),
                ("11111011000111001110111100110011001110011011010011010000100011011110110000100001101111011110111101110000101000101111011110111010000100001001010010100001000010011101011010100110110001100110011100111111"),
                ("11111111111111011110111100110010011100110100101001010000100011011110111011110111010000100001000101110000100001000010000111011010000100101001010010100101001010011001110011101101111001110111111111111111"),
                ("11111111111111011110011001100101001010010100001000010011100001000010001101101000110111011110111101110000100001000010000111011010000100001000010000100001000010011001110011101100110011110111111111111111"),
                ("11111111110111001110111011001111000110000100001000010010100101000010000100010111101111011110111000010000110111000010000111011010000100001000010000100001000010001100011000100111001111110111101111011111"),
                ("11111111110110001100110011001101000010000100001000010000100011011110111101110111000010000100001000011011110111000010000100001101110100001000010000100001000010000100101001110101011011001011000110001100"),
                ("11111111110110001100110011001101000010000100001000010000100011011110111101110111000010000100001000011011110111000010000100001101110100001000010000100001000010000100101001110101011011001011000110001100"),
                ("11111111111011010110101101001101001010010100001000010000100001000010001101100001000010000100001101111101111011010000100001000101111011111011110110100001000010000100001000110101011010011110011100111001"),
                ("11111111111011010110101101011011010110100100001000010000100001000010000100010111101111011110111101110000110111010000100010111000010000100001000011101101000010000100001000110101011010011110011100111001"),
                ("01110011001011010110100111001111010110100100101000010000100001001010010100011011101111011110111000010000100001101111011110111000011101101000010000100001000010000100001000100111001101100111101111011110"),
                ("01100111101001110011110101100001001010010100001001010010100001001010010100010111000010000100001000010000110111110111101110111010000100001000010000100001000010000100101001101101100111110111101111011111"),
                ("01100111101001110011110101100001001010010100001001010010100001001010010100010111000010000100001000010000110111110111101110111010000100001000010000100001000010000100101001101101100111110111101111011111"),
                ("11001011001100111001100110100111000110000100001001010010100011000110000100110111101110000100001000010000100001101111011111011010000100001000010000100001000010000100001000100111100111110111111111111111"),
                ("11001110011100111001100111101010011100110100101000010011100001001010010100011011010001011110111000010000100001000010000100001110110100001000010000100001001010010100101001100110110001110111111111111111"),
                ("11001110011001110011100111011010011100110100101000010000100101000010000100001000010001011110111000010000100001000010000110111010000100001000010000100001000110101001110011100110110011110111111111111111"),
                ("11111110011001110011101101001111000110000100101000010000100001000010000100001000010001101111011101110000100001000010000100001101110100001000010000100001000110101011010110101100110001110111111111111111"),
                ("11111110011001110011101101001111000110000100101000010000100001000010000100001000010001101111011101110000100001000010000100001101110100001000010000100001000110101011010110101100110001110111111111111111"),
                ("11111111111101011010100111101001001010011101001000010000100001000010000100001000010000100001000101111011100001000010000110111010000100001000010000100001000100111011010110101100110001110111111111111111"),

                -- explosion_3-4.png
                ("11111111110111001110011001011010110101101001101000010000100001000010000100010111000010000100001101111011101000010000100001000010000100001000010000100001000110100100101001110101001111010111111111111111"),
                ("11111111110111001110011001011010110101101101001000010000100001000010001011100001000010000100001000011011111011010000100001000010000100001000010000100001000010011100011000100111011010011110011100111111"),
                ("11111111111111011110011001001110011100111101001000010000100001000010000100010111000010000100001000010000110111010000100001000010000100001001010010100001000010011001110011101101001110011110011100111001"),
                ("11111111111111011110011001001110011100111101001000010000100001000010000100010111000010000100001000010000110111010000100001000010000100001001010010100001000010011001110011101101001110011110011100111001"),
                ("11111111110111001110011001001101001010010100101001010000100001000010001101100001000010000100001000010000110111010000100011011010000100111000110000100101000010011001110011110101001111001110011100111001"),
                ("11111111111111011110110011001101000010000100001000010000100001000010000100011011101110000100001000010000100001101111011110111010011100001000010000100101001010001100011000010011001111001011000110011001"),
                ("11111111101111011110110011011001001010010100001000010000100001000010000100010111110111011110111000010000100001000010000110111010000100101000010000100101001010000100101001110001101010011111101111001100"),
                ("11111111101111011110110011011001001010010100001000010000100001000010000100010111110111011110111000010000100001000010000110111010000100101000010000100101001010000100101001110001101010011111101111001100"),
                ("11110111100110001100100111001101000010000100001000010000100011011110110000110111101110000100001000010000110111101111011111011010000100101000010000100001000010011101011010100111001110110011000110001110"),
                ("11001110011001110011101101101001000010000100001000110110000100001000010000110111010001011110111000011011110111101111011110111010000100001000010000100001000010001101011010101101011010110111111111111111"),
                ("11001110011001110011101101101001000010000100001000010001101110111101111011101000010001101111011110111011100001000010000100001110110100001000010000100001000010000100101001100111011010110111111111111111"),
                ("01100011001100111001101101101001001010010100001000010000100001000010001011100001000011011110111101110000100001000010000110111110111101101000010000100001000010000100001000100111100101100111111111111111"),
                ("11111111101111011110100111001111000110000100001000010000100001000010000100011011000011011110111000010000110111101111011110111010000100001001010010100101000010001100011000100111110101110111111111111111"),
                ("11111111101111011110100111001111000110000100001000010000100001000010000100011011000011011110111000010000110111101111011110111010000100001001010010100101000010001100011000100111110101110111111111111111"),
                ("11111111111111011110011001011010011100110100101000010000100001000010000100011011000010000100001000011011110111110111101101000110110100011000110000100101000010000100101001110010110011110111111111111111"),
                ("11111111110111001110111101011010011100110100101001010010100101001010010100011011000010000100001000011011101000010000100010111101111101101000010000100001001010011001110011011001111011110111111111111111"),
                ("11111110010110001100011001001111010110100100101000010000100101000010000100010111101110100001000000011011110111101111011100001000011101101000010000100010011101101100111001011001111001110011000110011111"),
                ("11001110011001110011100111100001001010010100001000010000100001000010000100011011000011101111011110111011100001101111011100001110110100001000010000100011010101101100111001110011111011110011000110011001"),
                ("11001110011001110011100111100001001010010100001000010000100001000010000100011011000011101111011110111011100001101111011100001110110100001000010000100011010101101100111001110011111011110011000110011001"),
                ("11001110011001110011110100100101001010010100001000010000100001000010000100001000101110000100001101111011110111000010000110111010000100001000010000100011010101101011010110100111001111001110011100111001"),
                ("11001110011101011010110100100101001010010100001000010000100001000010000100001000101111011110111000010000110111000010000110111010000100001001010010100111010101101011010110101100110011001110011100111110"),
                ("01100011001001110011100111101011010110101100001000010000100001000010000100001000110111011110111010000100011011101111011110111010000100001000010000100101001110001001110011101101011011101011000110011110"),
                ("11111111011100111001101101011010110101101011011010010000100001000010000100001000110111101111011010000100001000010000100001000010000100001000010000100001001010011101011010101101001111110111101111011111"),
                ("11111111011100111001101101011010110101101011011010010000100001000010000100001000110111101111011010000100001000010000100001000010000100001000010000100001001010011101011010101101001111110111101111011111"),
                ("11111111111100111001101101011010110101101011011010010010100001000010000100001000110110100001000010000100001000010000100001000010000100101001010010100001000010011101011010101101100111101111111111111111"),
                ("11111111110110001100110011100110110101101011011010010010100001000010000100001000010000100001000010000100001000010000100001000010010100101000010000100001001010011101011010100111100111110111111111111111"),
                ("11111111110110001100011001100110011100111011010011010000100101001010010100001000010000100001000010000100101000010000100001000010010100101001010010100001000010010100101001110101100101100111111111111111"),
                ("11111111111100111001101101011010110101101001101001010010100101000010000100001000010000100001000010000100101001010010100101000010000100101001010010100001001010010100101001110001001110011111111111111111"),
                ("11111111111100111001101101011010110101101001101001010010100101000010000100001000010000100001000010000100101001010010100101000010000100101001010010100001001010010100101001110001001110011111111111111111"),
                ("11111111110110001100101101011011001110011101001001110000100101001010010100101000010000100001000010010100111010110001100001001010000100001000010000100001001110000100101001110101011011001111111111111111"),
                ("11111111111111111111101101111001100011001001110011110000100111010110101011010011010010100101001010011100010011110001100001001010010100001000010000100001000110000100101001110101011011111111111111111111"),
                ("11111111111111111111111110111011001110011100110110110100100111010110101011010110110000100101001110001001110110100111001101001110000100111000110000100111010110100100101001110101111111111111111111111111"),
                ("11111111111111111111111111111101100011000110010110100111100010011100111011010011110101101011010110101011010011100111001110110100111101001001010010100110011100111101011010100111111111111111111111111111"),
                ("11111111111111111111111111111101100011000110010110100111100010011100111011010011110101101011010110101011010011100111001110110100111101001001010010100110011100111101011010100111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111001100101101101011010110101011010011101101011010110100111011010011100111001110110101101101001001010011101010011101101011010110101101111111111111111111111111"),
                ("11111111111111111111111111111111111111111111110011100111001110110101101001110011100111011010110101101011010110101101011010110101101001110011100111011010110101101011010110111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111011000110011001110011100111001100111011010110101101011010110101101011010110101101011011001110011100110110101101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111110110011010110101001110011100111100111001101101011010110100111001110011100111100111001110011111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111110110011010110101001110011100111100111001101101011010110100111001110011100111100111001110011111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111101001001010010100101001100111100111001100111001110011110011100111001110011100111101111011111111111111111111111111111111111111111111111111111001"),

                -- explosion_3-5.png
                ("11111111111100111001110011100101100011000111011111111111111111111111111111111111111111100111001110011111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001"),
                ("11111110011100111001110010110011110111100110011111111111111111111111111111111111011000110001100110011100101100111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11010100111001110011110011100110011100111011010110101100110001110011101111011110011101111011110110011100111101111101111011101111100110010011100111100111111111111111111111111111111111111111111111111111"),
                ("11010100111001110011110011100110011100111011010110101100110001110011101111011110011101111011110110011100111101111101111011101111100110010011100111100111111111111111111111111111111111111111111111111111"),
                ("10011101101001110011100111001111010110101001110110101101100111101111010110011110111101111011110100110110010110100111001111001110011100110011100111011010110111111111111111111111111111111111111111111111"),
                ("11010100111011010110110100100111000110001001110110100111001110011100111100101100011001100111001100111011010110101101011010110100111101011000110001101011010110101001110011101101111111111111111111111111"),
                ("01001110001001110011100111100001001010011101011010010010100011000110000100110011110011100111001101101011010011110101101011010110100100101001010010100101001010011101011010101101011011111111111111111111"),
                ("01001110001001110011100111100001001010011101011010010010100011000110000100110011110011100111001101101011010011110101101011010110100100101001010010100101001010011101011010101101011011111111111111111111"),
                ("11010010010100101001010010100001000010000100101000010000100001000010000100001001101101011010110101101011011000010010100101001010010100101001010011100011000110101001110011101101011010110111111111111111"),
                ("01000010000100001000010000100101001010010100001000010000100001000010000100001001100111101011010110101101001001010010100101000010010100001001010010100101000110101001110011100111011010110111111111111111"),
                ("01000010000100001000010010100101001010010100001000010000100001001010010100101000010000100001000010000100101001010000100001000010000100001000010000100001000010010100101001110101011011001111111111111111"),
                ("01000010000100101001110000100001000010000100001000010000100001001010011100001000010000100001000010000100101000010000100001001010000100101001010010100001000110000100101001010011001111001110011100111101"),
                ("01000010000100001000010011100001001010010100101000010001101101000010000100011011110110100001000010000100001000010000100001001010010100101001010010100001000010011101011010110101001110110110011100111001"),
                ("01000010000100001000010011100001001010010100101000010001101101000010000100011011110110100001000010000100001000010000100001001010010100101001010010100001000010011101011010110101001110110110011100111001"),
                ("01000010000100001000010000100101000010000100001000110111101101000010001101110111000011101111011010000100001000010000100001000010010100101000010000100001001110001001110011101101011010110100111001111001"),
                ("01000010000100001000110111011110111101111101110111000011011110111101110100010111000010000100001101111011110111010000100001000010000100001000010000100101001010011011010110101101011010110100111001111001"),
                ("01000010000100001000010001011100001000011011110111000010000110111101111101101000101111011110111000010000110111010000100001000010000100001001010011100011000100111001110011100111011010110100111001111001"),
                ("01000110111011110111101110000100001000011011110111000010000110111101111011101000101110000100001101111011111011010000100001000010000100001001010011101010011101101001110011100111011010110101101011010011"),
                ("01000110111011110111101110000100001000011011110111000010000110111101111011101000101110000100001101111011111011010000100001000010000100001001010011101010011101101001110011100111011010110101101011010011"),
                ("10111101110000100001000010000100001000010000110111101110000100001000011011110111101111011110111101110000101000010000100001000010000100101001010010100111000100111011010110101101011010110101101011010011"),
                ("10111000010000100001000010000100001000010000100001110111011100001000010000100001000011101111011101110000101000010000100001000010000100001000010000100101001110001101011010100111011010110101101011010011"),
                ("00001000010000100001000010000110111101110000110111110111011110111101110000100001010001101111011000011011110111110111101101000010000100001000010000100001001010011101011010101101011010110110011100111001"),
                ("00001000010000100001000011011111011110111011101000010000000100001000010000100001101110000100001101111011111011110111101111011010000100001000010000100001001110001101011010101101001110011100111001110011"),
                ("00001000010000100001000011011111011110111011101000010000000100001000010000100001101110000100001101111011111011110111101111011010000100001000010000100001001110001101011010101101001110011100111001110011"),
                ("10111000011011110111000011101110111101111011110111010000000111011110111101111011101111101111011010000100001000010000100001000010000100001000010000100010011101101001110011100111001111001100111001101001"),
                ("01000101110100001000110110100001000010000000100001101111011101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100110110101101011010110101101001111001100111001101001"),
                ("01000010000100001000010000100001000010001101100001101110100001000010000100001001010000100001000010000100001000010000100001000010000100101000010000100111010110101001110011110101011011001110101101001001"),
                ("01000010000100001000010000100001000010000100000001110110100001000010000100001001010010100001000010000100001000010000100001000010000100101001010010100101001010011100011000110101001101100011000110011010"),
                ("01000010000100001000010000100001000010000100000001110110100001000010000100001001010010100001000010000100001000010000100001000010000100101001010010100101001010011100011000110101001101100011000110011010"),
                ("01000010000100001000010000100001000010000100011011010000100001000010000100001001010000100001000010000100001000010000100001001010010100001001010011100011000110101001110011101101001101100111111111111111"),
                ("01000010000100001000010010100001000010000100001000010000100001000010000100001001010000100001000010000100001000110101101011010110101001101001010010100110011101101011010110011001001111111111111111111111"),
                ("10011110101101011010010010100001000010000100001000010000100001000010000100101001010010100001000010000100011000101101011010110101101011010011100111101010011110010110001100111101111111111111111111111111"),
                ("10110101101001110011010010100001001010010100001000010000100111000110001001110011110100100101001010010100111010101101011010110101101001110110101101100101100110010110001100111111111111111111111111111111"),
                ("10110101101001110011010010100001001010010100001000010000100111000110001001110011110100100101001010010100111010101101011010110101101001110110101101100101100110010110001100111111111111111111111111111111"),
                ("10110101101001110011100111001110110101101001111010110101101010011100111011010110100111100011000010010100111010101101011010110110011100110110101101011011110011101111111111111111111111111111111111111111"),
                ("01100011000110001100011001100111001110011001110110101101011010011100110110011110011001001110011110101101010011101101011010110110010110010110101101011010110111111111111111111111111111111111111111111111"),
                ("01110011101111011110011101111011110111100110010011100111100111110111101111001110011001001110011100111101010011110011100111001011000110011001110010110011111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111110111101111011001110010110011110111101111111111110011100111001110011100101100111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111110111101111011001110010110011110111101111111111110011100111001110011100101100111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111011001110010110011111111111111111111111111100111001110011100101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- explosion_3-6.png
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001100110011100111001111111111111111111111111101100011001100111001111101111111111111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111010110001100110011100111001110011100111111111111111001100011001100111001111101111011110111111111111111111111111111111"),
                ("11111111111111111111111111111111111111111111111111011001100101100011000110011001110011001110011110101001110011011000110001110111101111011001110011001110011011001111011110111100111011110011100111001110"),
                ("11111111111111111111111111111111111111111111111111011001100101100011000110011001110011001110011110101001110011011000110001110111101111011001110011001110011011001111011110111100111011110011100111001110"),
                ("11111111111111111111111111111111111111111111110110101101011001100011001100110110101101001110011110101101010011011000110011110011001001110110101101011010110100111100111001110010110001100011000110001100"),
                ("11111111111111111111111111111111111111110111011110101101011011001110011100110110101101101011010010010100111000100111001110110101101001111010110101101011010100111011010110100111001110011101101011010110"),
                ("11111111111111111111111111111101100011001100101100110011011010011100111011010110101101101011010010010100101001110101101010011100111100001001010010100001000010000100101001010000100110011101101011010110"),
                ("11111111111111111111111111111101100011001100101100110011011010011100111011010110101101101011010010010100101001110101101010011100111100001001010010100001000010000100101001010000100110011101101011010110"),
                ("11111111111111111111111111111001100011001100110011110101001110110101101011010110101101100011000010000100001000010010100101001010010100001000010000100001000010000100001000010000100111010110101101010011"),
                ("11111111111111111111100110110010110101101011010011010010100110011100111101011010110100100001000010000100001000010000100001001010000100001000010000100001000010000100001000010000100101000010000100001000"),
                ("11111111110110001100100111011010011100111101011000110000100101000010000100101001010000100001000010000100001000010000100001001010000100001000010000100011011010000100001000010000100001000010000100001000"),
                ("11010011000110001100100111101011000110000100101001010010100101001010010100001000010000100001000010000100001000010010100101001010000100001000010001101100001010000100001000010000100001000010000100001000"),
                ("01001110101100111001101101101010011100111101011010010010100001001010010100001000010000100001000010000100001000010000100001001010000100001000010001011100001110110100001000010000100001000010000100001000"),
                ("01001110101100111001101101101010011100111101011010010010100001001010010100001000010000100001000010000100001000010000100001001010000100001000010001011100001110110100001000010000100001000010000100001000"),
                ("01001100111100111001100111011010110101101011010110010010100001000010000100001000010000100001000010000100001000010000100001000010000100010111101111011100001000010100001000010001101101000101111011101000"),
                ("01001100111100111001100111001110011100111011010011010000100001000010000100001000010000100001000010000100011011101111011111011110111101100001000010100010111101111011110111110110000110111000010000110111"),
                ("10011100111001110011100111011011010110101100001001010000100001000010000100011011110111101111011101111011100001101111011100001000010000100001000010100001000101111101111011101110000100001000010000100001"),
                ("11001110011011010110101101011011010110100100101001010000100001000010000100001000110111011110111101110000111011010000100000001000011011110111101111101110111000011011110111000010000100001000010000100001"),
                ("11001110011011010110101101011011010110100100101001010000100001000010000100001000110111011110111101110000111011010000100000001000011011110111101111101110111000011011110111000010000100001000010000100001"),
                ("10011101101011010110101101001111010110101100001001010010100001000010000100001000010000100001000000011011111011000010000100001000010000110111101111101100001000010000100001000010000100001000010000110111"),
                ("10011101101011010110101101011010110101101001111000010010100101001010010100001000010000100001000000011011110111101111011110111101110000100001000011011110111000010000100001000010000100001101111011110111"),
                ("10011101101011010110101101001110011100111011010011110100100101000010000100001000010001101111011101111011100001101111011101000101111011100001000010000110111101110000100001000011011110111110111101101000"),
                ("11001100111011010110101101001110011100111001111000110000100101000010000100001000010001011110111000010000110111101111011101000110111011100001000010000110111101110000100001101110100001000010000100001000"),
                ("11001100111011010110101101001110011100111001111000110000100101000010000100001000010001011110111000010000110111101111011101000110111011100001000010000110111101110000100001101110100001000010000100001000"),
                ("11001100111011010110101101011010110101100100101001010010100001000010000100001000010001011110111101111011100001000010000110111010001011110111101110000110111110111011110111101111101101000010000100001000"),
                ("11001100111011010110101101011010011100111100001001010000100001001010010100101000010000100001000010000100011011000010000110111110110100011011110111101101000010000100001000010010100001000010000100001000"),
                ("11001110011011010110100111101011010110100100101000010000100101001010010100101001010000100001000010000100001000110111101111011010000100011011110110100001000010010100101001110000100101000010000100001000"),
                ("11101110011100111001100110100101001010011100001000010000100101001010010100001001010000100001000010010100001000010000100001000110000100101000010000100001000010000100001000010001100001001010000100001000"),
                ("11101110011100111001100110100101001010011100001000010000100101001010010100001001010000100001000010010100001000010000100001000110000100101000010000100001000010000100001000010001100001001010000100001000"),
                ("11111111111100111001101101101001001010010100101000010000100001000010000100001000010000100101001010010100001000010000100001000010010100101000010000100001000010000100101001010010100101000010000100001000"),
                ("11111111111011010110101101001110011100111101001000010010100101000010000100101000010010100101001110101101011010100111001101001010000100001000010000100001000010000100101001010010100001000010000100001000"),
                ("11111111111011010110101101011010011100111101011000110000100101001010010100101001010011100011000101101011010110101101011001001010000100001000010000100001000010010100001000010000100101001010010100111010"),
                ("11111111111111111111101101011011010110100100101001010010100101001010011101011010110101001110011101101011011001110011100110011010011100001000010000100111010110100100101001110001001110011110001100001001"),
                ("11111111111111111111101101011011010110100100101001010010100101001010011101011010110101001110011101101011011001110011100110011010011100001000010000100111010110100100101001110001001110011110001100001001"),
                ("11111111111111111111111111011010011100111101011010110101100011010110101001110110101101011010110101101001111001011000110001100110011001110011100111001110110100111100011000010011101010110100111001111010"),
                ("11111111111111111111111111111111111111111111110110101101001111001110011100111001100111011010110011001001111110111101111011110011001110111001110011011010110100111101011010100111001110011101101011010011"),
                ("11111111111111111111111111111111111111111111111111110011001101100011001111011101111101110111101110011100111110011100111011110111100111001100011001011010110101101001110011110011100110011100111001111010"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001100110011100101100011000110011111111111111111111111111111111111011001111011110011001100111001110011100111111"),
                ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111100110001100110011100101100011000110011111111111111111111111111111111111011001111011110011001100111001110011100111111"),
                ("11001111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111101100111001111111111111111111111111111111111111111111111011100110001100110011100111001111111111111111"),

                -- unbreakeable_1.bmp
                ("11101111010111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110010000100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100100001000001100011000110111101111"),
                ("11101111010111101111011110010000100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100100001000001100011000110111101111"),
                ("11101111010111101111011110010000100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100100001000001100011000110111101111"),
                ("11101111010111101111011110000100001000010000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110000100001000010000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010001100011000110111101111"),
                ("11101111010111101111011110000100001000010000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110000100001000010000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110000100001000010000100001001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010001100011000110111101111"),
                ("11101111010111101111011110010000100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100100001000001100011000110111101111"),
                ("11101111010111101111011110010000100000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100100001000001100011000110111101111"),
                ("11101111010111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110111101111"),
                ("11101111010111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110111101111"),
                ("11101111010111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110111101111"),
                ("11101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("11101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("11101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("11101111011110111101111011111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110"),
                ("11101111011110111101111011111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110"),
                ("11101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011111011110"),
                ("11101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011111011110"),
                ("11101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011111011110"),
                ("11100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100"),
                ("11100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100"),

                -- unbreakeable_2.bmp
                ("11100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("11100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("11100111000111101111011110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000001100011000111110111101"),
                ("11100111000111101111011110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000001100011000111110111101"),
                ("11100111000111101111011110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000001100011000111110111101"),
                ("11100111001111011110111100001100011000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100001100011000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011001000010000100001000010000011000110001100011001000010000100001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011001000010000100001000010000011000110001100011001000010000100001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011001000010000100001000010000011000110001100011001000010000100001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011011110111100100001000010000011000110001100011011110111101111001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011011110111100100001000010000011000110001100011011110111101111001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011001000010000100001000010000011000110001100011001000010000100001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011001000010000100001000010000011000110001100011001000010000100001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011011110111100100001000010000011000110001100011011110111101111001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011011110111100100001000010000011000110001100011011110111101111001000010001111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110111101111011111110111101"),
                ("11100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011111110111101"),
                ("11100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011111110111101"),
                ("11100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011111110111101"),
                ("11100111001111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100111101111011111110111101"),
                ("11100111001111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100111101111011111110111101"),
                ("11100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("11100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("11100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("11100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110111101"),
                ("11100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110111101")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 2515 := 0;
    out_color_reg : std_logic_vector(4 downto 0) := (others => '0');
begin
    process(in_sprite_nb, in_sprite_row, in_sprite_col)
    begin
        case in_sprite_nb is
            when 0 => real_row <= in_sprite_row;
            when 1 => real_row <= 40 + in_sprite_row;
            when 2 => real_row <= 107 + in_sprite_row;
            when 3 => real_row <= 174 + in_sprite_row;
            when 4 => real_row <= 241 + in_sprite_row;
            when 5 => real_row <= 281 + in_sprite_row;
            when 6 => real_row <= 321 + in_sprite_row;
            when 7 => real_row <= 361 + in_sprite_row;
            when 8 => real_row <= 401 + in_sprite_row;
            when 9 => real_row <= 462 + in_sprite_row;
            when 10 => real_row <= 523 + in_sprite_row;
            when 11 => real_row <= 584 + in_sprite_row;
            when 12 => real_row <= 645 + in_sprite_row;
            when 13 => real_row <= 706 + in_sprite_row;
            when 14 => real_row <= 767 + in_sprite_row;
            when 15 => real_row <= 828 + in_sprite_row;
            when 16 => real_row <= 889 + in_sprite_row;
            when 17 => real_row <= 950 + in_sprite_row;
            when 18 => real_row <= 1011 + in_sprite_row;
            when 19 => real_row <= 1072 + in_sprite_row;
            when 20 => real_row <= 1133 + in_sprite_row;
            when 21 => real_row <= 1194 + in_sprite_row;
            when 22 => real_row <= 1255 + in_sprite_row;
            when 23 => real_row <= 1316 + in_sprite_row;
            when 24 => real_row <= 1356 + in_sprite_row;
            when 25 => real_row <= 1396 + in_sprite_row;
            when 26 => real_row <= 1436 + in_sprite_row;
            when 27 => real_row <= 1476 + in_sprite_row;
            when 28 => real_row <= 1516 + in_sprite_row;
            when 29 => real_row <= 1556 + in_sprite_row;
            when 30 => real_row <= 1596 + in_sprite_row;
            when 31 => real_row <= 1636 + in_sprite_row;
            when 32 => real_row <= 1676 + in_sprite_row;
            when 33 => real_row <= 1716 + in_sprite_row;
            when 34 => real_row <= 1756 + in_sprite_row;
            when 35 => real_row <= 1796 + in_sprite_row;
            when 36 => real_row <= 1836 + in_sprite_row;
            when 37 => real_row <= 1876 + in_sprite_row;
            when 38 => real_row <= 1916 + in_sprite_row;
            when 39 => real_row <= 1956 + in_sprite_row;
            when 40 => real_row <= 1996 + in_sprite_row;
            when 41 => real_row <= 2036 + in_sprite_row;
            when 42 => real_row <= 2076 + in_sprite_row;
            when 43 => real_row <= 2116 + in_sprite_row;
            when 44 => real_row <= 2156 + in_sprite_row;
            when 45 => real_row <= 2196 + in_sprite_row;
            when 46 => real_row <= 2236 + in_sprite_row;
            when 47 => real_row <= 2276 + in_sprite_row;
            when 48 => real_row <= 2316 + in_sprite_row;
            when 49 => real_row <= 2356 + in_sprite_row;
            when 50 => real_row <= 2396 + in_sprite_row;
            when 51 => real_row <= 2436 + in_sprite_row;
            when 52 => real_row <= 2476 + in_sprite_row;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= (rom(real_row))(((in_sprite_col + 1) * 5 - 1) downto (in_sprite_col * 5));
        end if;
    end process;
    out_color <= out_color_reg;
end behavioural;
