


entity collision_detector_rect_rect
port(
    x : vector;
    width, height : 
);
end game_controller;


architecture behavioural of game_controller is

-- Choices

begin


-- Map generation

end architecture;
