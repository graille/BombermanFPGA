library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.PROJECT_PARAMS_PKG.all;
use work.PROJECT_TYPES_PKG.all;
use work.PROJECT_DIRECTION_PKG.all;

entity font_sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_id : in block_category_type;
        in_sprite_state : in state_type;
        in_sprite_direction : in direction_type;

        in_sprite_row : in integer range 0 to 36;
        in_sprite_col : in integer range 0 to 27;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end font_sprite_rom;

architecture behavioral of font_sprite_rom is
    subtype word_t is std_logic_vector(0 to 139);
    type memory_t is array(0 to 3551) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- 0_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 1_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 2_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff8000003fff800007ffffffff"),
                (x"fffffffffff8000003ff0000007ffffffff"),
                (x"fffffffffff8000003ff0000007ffffffff"),
                (x"fffffffffff8000003ff0000007ffffffff"),
                (x"fffffffffff8000003ff0000007ffffffff"),
                (x"fffffffffff8000003e00000007ffffffff"),
                (x"fffffffffff8000003e000000ffffffffff"),
                (x"fffffffffff8000003e000000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 3_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffe00000007ffffffff"),
                (x"ffffffffe000000fffe00000007ffffffff"),
                (x"ffffffffe000000fffe00000007ffffffff"),
                (x"ffffffffe000000fffe000000ffffffffff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffffffffe000000fffff00000ffffffffff"),
                (x"ffffffffe00000007fff00000ffffffffff"),
                (x"ffffffffe00000007fff00000ffffffffff"),
                (x"ffffffffe00000007fff00000ffffffffff"),
                (x"ffffffffff0000007fff00000ffffffffff"),
                (x"ffffffffff00000fffff00000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 4_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffff8000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff0000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffe0000000000000000003fffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe000000f800007fffffffffffff"),
                (x"ffffffffe000000f800007fffffffffffff"),
                (x"ffffffffe000000f800007fffffffffffff"),
                (x"ffffffffe000000f800007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"fffffffffff80000000000000003fffffff"),
                (x"ffffffffffffffff800000000003fffffff"),
                (x"ffffffffffffffff8000000000001ffffff"),
                (x"ffffffffffffffff8000000000001ffffff"),
                (x"ffffffffffffffff800007fe00001ffffff"),
                (x"ffffffffffffffff800007fe00001ffffff"),
                (x"ffffffffffffffff800007fe00001ffffff"),
                (x"ffffffffffffffff800007fe00001ffffff"),
                (x"ffffffffffffffff8000000000001ffffff"),
                (x"ffffffffe00000000000000000001ffffff"),
                (x"ffffffffe0000000000000000003fffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 5_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff80000000007ffffffffffffffffff"),
                (x"fffe0000000000007ffffffffffc00003ff"),
                (x"fffe0000000000007ffffffff000000001f"),
                (x"fffe00000000000003fffffe0000000001f"),
                (x"fffe00000000000003fff800000000003ff"),
                (x"fffe00000000000003ff0000000000003ff"),
                (x"fffe00000000000003ff0000000000003ff"),
                (x"ffffff80000000007fff00000003fffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffff800000000000000001ffffff"),
                (x"ffffffffff00000003e0000000001ffffff"),
                (x"ffffffffff00000003e0000000001ffffff"),
                (x"ffffffffe00000007fe0000000001ffffff"),
                (x"ffffffffe00000007fe0000000001ffffff"),
                (x"ffffffffe00000007fe0000000001ffffff"),
                (x"ffffffffe000000fffe0000000001ffffff"),
                (x"ffffffffe000000fffff00000003fffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 6_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 7_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 8_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"fffffffc0007fffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"fffffffffffffff0000000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 9_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc000000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"fffffffffffffffffc000000007ffffffff"),
                (x"fffffffffffffffffc000000007ffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff8000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 10_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffffffffff8000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 11_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000000000001ffffff"),
                (x"fffffffffffffff00000000000001ffffff"),
                (x"fffe0000000000000000000000001ffffff"),
                (x"fffe0000000000000000000000001ffffff"),
                (x"fffe0000000000000000000000001ffffff"),
                (x"fffe00000000000000000001fffffffffff"),
                (x"fffe0000000000000000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 12_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 13_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"f80000000000000000000000000000fffff"),
                (x"f80000000000000000000000000000fffff"),
                (x"f80000000000000000000000000000fffff"),
                (x"f80000000000000000000000000000fffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 14_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 15_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 16_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc0000000fffe00001ffffff"),
                (x"fffffffffff800000000000000001ffffff"),
                (x"ffffffffe00000000000000000001ffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"ffffff8000003fffffe00000007ffffffff"),
                (x"ffffff8000003fffffe00000007ffffffff"),
                (x"ffffff8000003ffffc000000007ffffffff"),
                (x"ffffff800007fffffc000000007ffffffff"),
                (x"ffffff800007ffff800000000003fffffff"),
                (x"ffffff800007fff0000000000003fffffff"),
                (x"ffffff800007fff0000000000003fffffff"),
                (x"ffffff800007c0000000f8000003fffffff"),
                (x"ffffff800007c0000000f8000003fffffff"),
                (x"ffffff800007c0000000f8000003fffffff"),
                (x"ffffff8000000000001ff8000003fffffff"),
                (x"ffffff800000000003fff8000003fffffff"),
                (x"ffffff800000000003fff8000003fffffff"),
                (x"ffffff80000000007ffff8000003fffffff"),
                (x"fffffffc000000007ffff8000003fffffff"),
                (x"fffffffc0000000fffff00000003fffffff"),
                (x"fffffffc0000000fffff00000003fffffff"),
                (x"ffffff800000000003e000000003fffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff800007c000000000000ffffffffff"),
                (x"fffffffffffffffffc0007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 17_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 18_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"fffe00000000000003fffffffffffffffff"),
                (x"fffe000000000000001ffffffffffffffff"),
                (x"fffe000000000000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 19_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc000000000000fffffffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffff80000000007ffffffff"),
                (x"ffffffffffffffff80000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff00000ffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 20_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffff800007ffffffff"),
                (x"fffffffc0000000ffffff800007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000000000fffff"),
                (x"ffffffffe000000000000000000000fffff"),
                (x"ffffffffe000000000000000000000fffff"),
                (x"ffffffffe000000000000000000000fffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 21_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"ffffff8000000000001ffffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"ffffffffffffffff800000000ffffffffff"),
                (x"fffffffffffffffffc000000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"fffffffffffffffffc0000000003fffffff"),
                (x"fffffffffffffffffc0000000003fffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 22_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe0003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc000000000000fffffffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc000000007c000000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffff00000003fffffff"),
                (x"fffffffc00003ffffffff8000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 23_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"ffffffffffffffff800000000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"ffffffffffffffff800000000ffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffff0000007ffffffffffffffffff"),
                (x"ffffffffff0000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 24_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc0000000ffc0000000ffffffffff"),
                (x"ffffff8000003fffffe000000ffffffffff"),
                (x"ffffff8000003fffffe000000ffffffffff"),
                (x"ffffff800007ffffffe000000ffffffffff"),
                (x"ffffff800007ffffffe000000ffffffffff"),
                (x"ffffff800007ffffffe000000ffffffffff"),
                (x"ffffff800007fffffc0000000ffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffc0000000003e00000007ffffffff"),
                (x"fffffffc0000000fffff0000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003ff000000000007ffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 25_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff0000007fe00000007ffffffff"),
                (x"ffffffffff0000007fe00000007ffffffff"),
                (x"ffffffffff0000007fe00000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 26_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 27_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 28_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"ffffffffffffffffffff000000001ffffff"),
                (x"ffffffffffffffffffff000000001ffffff"),
                (x"ffffffffffffffffffe0000000001ffffff"),
                (x"ffffffffffffffff8000000000001ffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"fffe00000000000003fffffffffffffffff"),
                (x"fffe0000000000007ffffffffffffffffff"),
                (x"fffe0000000000007ffffffffffffffffff"),
                (x"fffe000000000000001ffffffffffffffff"),
                (x"fffe000000000000001ffffffffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffffffc000000000000003fffffff"),
                (x"ffffffffffffffff8000000000001ffffff"),
                (x"fffffffffffffffffc00000000001ffffff"),
                (x"fffffffffffffffffc00000000001ffffff"),
                (x"fffffffffffffffffffff80000001ffffff"),
                (x"fffffffffffffffffffffffff0001ffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 29_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe00000007fffffffffffffffffffffff"),
                (x"fffe00000000000000000000007ffffffff"),
                (x"fffe00000000000000000000007ffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 30_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"fffe00000000000ffffffffffffffffffff"),
                (x"fffe00000000000003fffffffffffffffff"),
                (x"fffe00000000000003fffffffffffffffff"),
                (x"fffe000000000000001ffffffffffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffffff800000000000000001ffffff"),
                (x"fffffffffffffff00000000000001ffffff"),
                (x"ffffffffffffffff80000000000000fffff"),
                (x"ffffffffffffffffffff0000000000fffff"),
                (x"ffffffffffffffff80000000000000fffff"),
                (x"ffffffffffffffff80000000000000fffff"),
                (x"ffffffffffffffff80000000000000fffff"),
                (x"ffffffffffffc00000000000007ffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"fffffffc00000000001ffffffffffffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0007fffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 31_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 32_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffff8000003ffffc000000007ffffffff"),
                (x"ffc000000007ffffffff00000003fffffff"),
                (x"ffc0000000000000001ff8000003fffffff"),
                (x"ffc000001ff80000000007fe0003fffffff"),
                (x"f8000003ff000000000007fe0003fffffff"),
                (x"f8000003ff000000000007fe0003fffffff"),
                (x"f8000003ff000000000000000003fffffff"),
                (x"f8000003ff000000000000000003fffffff"),
                (x"f8000003ff000000000000000003fffffff"),
                (x"f8000003ff000000000000000003fffffff"),
                (x"f80000001f000000000000000003fffffff"),
                (x"f800000000000000000000000ffffffffff"),
                (x"ffc000000000000000000001fffffffffff"),
                (x"fffe000000003ffffffffffffffffffffff"),
                (x"fffe000000003ffffffffffffffffffffff"),
                (x"ffffff800000000003fffffe00001ffffff"),
                (x"fffffffc000000000000000000001ffffff"),
                (x"fffffffc000000000000000000001ffffff"),
                (x"ffffffffff0000000000000000001ffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 33_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffff8000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"fffffffc0000000f800007fffffffffffff"),
                (x"fffffffc00003fff800007fffffffffffff"),
                (x"fffffffc00003fff800007fffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff800007ffff80000001fffffffffff"),
                (x"fffe00000007fffffc000001fffffffffff"),
                (x"fffe000000fffffffc000000007ffffffff"),
                (x"fffe000000fffffffc000000007ffffffff"),
                (x"fffe000000fffffffc000000007ffffffff"),
                (x"fffe000000ffffffffe00000007ffffffff"),
                (x"fffe000000ffffffffff0000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 34_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"fffe000000000000000007fffffffffffff"),
                (x"fffe000000ffffff80000001fffffffffff"),
                (x"fffe000000ffffff80000001fffffffffff"),
                (x"fffe000000ffffff80000001fffffffffff"),
                (x"fffe000000fffffffc000001fffffffffff"),
                (x"fffe000000ffc00000000001fffffffffff"),
                (x"fffe000000f8000000000001fffffffffff"),
                (x"fffe00000000000000000001fffffffffff"),
                (x"fffe000000000000000007fffffffffffff"),
                (x"fffe00000000000000000001fffffffffff"),
                (x"fffe00000000000000000001fffffffffff"),
                (x"fffe000000003fff800000000ffffffffff"),
                (x"fffe000000fffffffc000000007ffffffff"),
                (x"fffe000000ffffffffff0000007ffffffff"),
                (x"fffe000000ffffffffff00000003fffffff"),
                (x"fffe000000ffffffffff00000003fffffff"),
                (x"fffe000000ffffffffe000000003fffffff"),
                (x"fffe000000ffffffffe000000003fffffff"),
                (x"fffe000000fffff000000000007ffffffff"),
                (x"fffe000000000000000000000ffffffffff"),
                (x"fffe00000000000000000001fffffffffff"),
                (x"fffe000000000000000007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 35_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff0000007fe00000007ffffffff"),
                (x"ffffffffe00000007fff0000007ffffffff"),
                (x"ffffffffe00000007fff0000007ffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffffffc00000000000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 36_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"fffffffc00000000001ffffffffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00003fff80000000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"ffffffffe0003fffffff0000007ffffffff"),
                (x"ffffffffe0003fffffff0000007ffffffff"),
                (x"ffffffffe0003ffffc000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 37_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe0003ffffffffffffffffffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00003ffffffffffe0003fffffff"),
                (x"fffffffc00003ffffffffffe0003fffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffff0000007ffffffffffffffffff"),
                (x"ffffffffff00000ffffffffffffffffffff"),
                (x"ffffffffff00000ffffffffffffffffffff"),
                (x"ffffffffff0000000000000000001ffffff"),
                (x"ffffffffff0000000000000000001ffffff"),
                (x"ffffffffff0000000000000000001ffffff"),
                (x"ffffffffff0000007fe0000000001ffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 38_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 39_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"fffffffffff80000000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffe00000007ffff800007ffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003fff8000000000001ffffff"),
                (x"fffffffc00003fff8000000000001ffffff"),
                (x"fffffffc00003fff8000000000001ffffff"),
                (x"fffffffc00003fff8000000000001ffffff"),
                (x"fffffffc00003fff8000000000001ffffff"),
                (x"ffffff8000003fffffff00000003fffffff"),
                (x"ffffff8000003ffffc0000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 40_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000fffffffffffffe00001ffffff"),
                (x"ffffff8000ffffffffff000000001ffffff"),
                (x"ffffff80000000000000000000001ffffff"),
                (x"ffffff80000000000000000000001ffffff"),
                (x"ffffff80000000000000000000001ffffff"),
                (x"ffffff80000000000000000000001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff8000003ffffffffffe00001ffffff"),
                (x"ffffff8000003ffffffffffe00001ffffff"),
                (x"ffffff8000003ffffffffffe00001ffffff"),
                (x"ffffff8000003ffffffffffe00001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 41_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 42_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc0000000000000001ffffff"),
                (x"ffffffffffffc0000000000000001ffffff"),
                (x"ffffffffffffc0000000000000001ffffff"),
                (x"ffffffffffffc0000000000000001ffffff"),
                (x"ffffffffffffc0000000000000001ffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc0000000fffe000000ffffffffff"),
                (x"fffffffc0000000ffc0000000ffffffffff"),
                (x"fffffffc0000000ffc0000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 43_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe0003ffffffffffffffffffffff"),
                (x"ffffffffe0003ffffffffffe0003fffffff"),
                (x"ffffffffe0003ffffffff8000003fffffff"),
                (x"ffffffffe0003fffffe000000003fffffff"),
                (x"ffffffffe0003fffffe000000003fffffff"),
                (x"ffffffffe0003fffffe000000003fffffff"),
                (x"ffffffffe0003ffffc0000000ffffffffff"),
                (x"ffffffffe0003fff80000001fffffffffff"),
                (x"ffffffffe0003ff0000007fffffffffffff"),
                (x"ffffffffe0003ff0000007fffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0003ff000000000007ffffffff"),
                (x"ffffffffe0003fff8000000000001ffffff"),
                (x"ffffffffe0003fffffe0000000001ffffff"),
                (x"ffffffffe0003fffffff0000000000fffff"),
                (x"ffffffffe0003fffffff0000000000fffff"),
                (x"ffffffffe0003ffffffffffe000000fffff"),
                (x"ffffffffe0003ffffffffffff00000fffff"),
                (x"ffffffffe0003fffffffffffff8000fffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 44_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffffffe0000000000000000003fffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 45_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe00000007ffffffffffffff8000fffff"),
                (x"fffe000000003ffffffffffff00000fffff"),
                (x"fffe00000000000ffffffffe000000fffff"),
                (x"fffe0000000000007ffffffe000000fffff"),
                (x"fffe000000000000001f0000000000fffff"),
                (x"fffe000000000000001f0000000000fffff"),
                (x"fffe00000000000000000000000000fffff"),
                (x"fffe000000f8000000000000000000fffff"),
                (x"fffe000000ffc00000000000000000fffff"),
                (x"fffe000000fffff000000001f00000fffff"),
                (x"fffe000000ffffff800007fff00000fffff"),
                (x"fffe000000fffffffc0007fff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 46_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe00001ffffffffffffffe00001ffffff"),
                (x"fffe00000007fffffffffffe00001ffffff"),
                (x"fffe000000003ffffffffffe00001ffffff"),
                (x"fffe00000000000ffffffffe00001ffffff"),
                (x"fffe00000000000ffffffffe00001ffffff"),
                (x"fffe00000000000ffffffffe00001ffffff"),
                (x"fffe0000000000007ffffffe00001ffffff"),
                (x"fffe00000000000003fffffe00001ffffff"),
                (x"fffe00001f000000001ffffe00001ffffff"),
                (x"fffe00001ff80000001ffffe00001ffffff"),
                (x"fffe00001fffc000001ffffff0001ffffff"),
                (x"fffe00001fffc0000000fffe00001ffffff"),
                (x"fffe00001ffffff0000007fe00001ffffff"),
                (x"fffe00001ffffff0000007fe00001ffffff"),
                (x"fffe00001ffffff00000000000001ffffff"),
                (x"fffe00001fffffff8000000000001ffffff"),
                (x"fffe00001ffffffffc00000000001ffffff"),
                (x"fffe00001fffffffffe0000000001ffffff"),
                (x"fffe00001ffffffffffff80000001ffffff"),
                (x"fffe00001ffffffffffff80000001ffffff"),
                (x"fffe00001ffffffffffff80000001ffffff"),
                (x"fffe00001ffffffffffff80000001ffffff"),
                (x"fffe00001ffffffffffffffffffffffffff"),
                (x"fffe00001ffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 47_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"ffffff800000000fffe000000003fffffff"),
                (x"ffffff800000000fffe000000003fffffff"),
                (x"fffe000000003ffffffff800000000fffff"),
                (x"fffe00000007fffffffffffe000000fffff"),
                (x"fffe000000fffffffffffffe000000003ff"),
                (x"fffe000000fffffffffffffff00000003ff"),
                (x"fffe000000ffffffffffffffff8000003ff"),
                (x"fffe000000ffffffffffffffff8000003ff"),
                (x"fffe000000ffffffffffffffff8000003ff"),
                (x"fffe000000ffffffffffffffff8000003ff"),
                (x"fffe000000ffffffffffffffff8000003ff"),
                (x"fffe000000ffffffffffffffff8000003ff"),
                (x"fffe00000007ffffffffffffff8000003ff"),
                (x"fffe000000003ffffffffffff00000003ff"),
                (x"ffffff80000000007ffffffff00000003ff"),
                (x"fffffffc0000000000000000000000fffff"),
                (x"fffffffc0000000000000000000000fffff"),
                (x"ffffffffe000000000000000000000fffff"),
                (x"ffffffffff0000000000000000001ffffff"),
                (x"ffffffffffffc000000000000003fffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 48_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc000000000000fffffffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0007ffff800000000003fffffff"),
                (x"fffffffc0007ffff800000000003fffffff"),
                (x"fffffffc0007ffffffe000000003fffffff"),
                (x"fffffffc00003ffffffff8000003fffffff"),
                (x"fffffffc00003ffffffff8000003fffffff"),
                (x"fffffffc00003fffffff00000003fffffff"),
                (x"fffffffc00003fffffe000000003fffffff"),
                (x"fffffffc00003ffffc000000007ffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"fffffffc00000000001ffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 49_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffe0000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00003ffffffff8000003fffffff"),
                (x"ffffff8000003ffffffff8000003fffffff"),
                (x"ffffff8000003ffffffff8000003fffffff"),
                (x"ffffff800007fffffffffffe0003fffffff"),
                (x"ffffff800007fffffffffffe0003fffffff"),
                (x"ffffff800007fffffffffffe0003fffffff"),
                (x"ffffff800007fffffffffffe0003fffffff"),
                (x"ffffff800007fffffffffffe0003fffffff"),
                (x"ffffff800007fffffc0000000003fffffff"),
                (x"ffffff800007fffffc0000000003fffffff"),
                (x"ffffff800007fffffc0000000003fffffff"),
                (x"ffffff800007fffffc0000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"ffffff8000000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"ffffffffe00000000000000000001ffffff"),
                (x"fffffffffffffffffffff80000001ffffff"),
                (x"fffffffffffffffffffffffe00001ffffff"),
                (x"fffffffffffffffffffffffe00001ffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 50_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"fffe00000000000000000001fffffffffff"),
                (x"fffe000000000000000000000ffffffffff"),
                (x"fffe00000007fffffc0000000ffffffffff"),
                (x"fffe00000007fffffc0000000ffffffffff"),
                (x"ffffff800007ffffffe000000ffffffffff"),
                (x"ffffff800007ffff80000001fffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff8000000000001ffffffffffffffff"),
                (x"ffffff8000000000001ffffffffffffffff"),
                (x"ffffff8000000000001ffffffffffffffff"),
                (x"ffffff8000000000001ffffffffffffffff"),
                (x"ffffff800007c000001ffffffffffffffff"),
                (x"ffffff800007c00000000001fffffffffff"),
                (x"ffffff800007c000000000000ffffffffff"),
                (x"ffffff800007ffff80000000007ffffffff"),
                (x"ffffff800007ffff80000000007ffffffff"),
                (x"ffffff800007ffff80000000007ffffffff"),
                (x"ffffff800007ffffffe00000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 51_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000000000000003fffffff"),
                (x"fffffffffff800000000000000001ffffff"),
                (x"ffffffffff0000000000000000001ffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"fffffffc000000007ffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"fffffffffffffffffc000000007ffffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"ffffffffffffffffffff00000003fffffff"),
                (x"fffffffffffffffffffff8000003fffffff"),
                (x"ffffffffff00000ffffff8000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 52_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe00000000000000000000007ffffffff"),
                (x"ffc000000000000000000000007ffffffff"),
                (x"ffc000000000000000000000007ffffffff"),
                (x"ffc000000000000000000000007ffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 53_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc0007fffffffffffffffffffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffff0001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc0007fffffffffffe00001ffffff"),
                (x"fffffffc00003ffffffffffe00001ffffff"),
                (x"fffffffc00003ffffffff80000001ffffff"),
                (x"fffffffc0000000ffffff80000001ffffff"),
                (x"fffffffc000000007fe000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 54_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffff00000fffff"),
                (x"fffe00001ffffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffe000000fffff"),
                (x"fffe00000007fffffffffffe000000fffff"),
                (x"fffe00000007fffffffffffe00001ffffff"),
                (x"ffffff800007fffffffff80000001ffffff"),
                (x"ffffff800007fffffffff80000001ffffff"),
                (x"ffffff800007fffffffff80000001ffffff"),
                (x"ffffff8000003ffffffff80000001ffffff"),
                (x"ffffff8000003ffffffff8000003fffffff"),
                (x"fffffffc0000000ffffff8000003fffffff"),
                (x"fffffffc000000007fe000000003fffffff"),
                (x"ffffffffe00000007fe00000007ffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 55_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffc00003fffffffffffffffffffffffffff"),
                (x"ffc00003ffffffffffffffffff8000fffff"),
                (x"ffc00003ffffffffffffffffff8000003ff"),
                (x"ffc00003fffffffffffffffff00000003ff"),
                (x"ffc00003fffffffffffffffff00000003ff"),
                (x"ffc00003fffffffffffffffff00000003ff"),
                (x"ffc000001ffffffffffffffff00000fffff"),
                (x"ffc000001ffffffffffffffff00000fffff"),
                (x"ffc0000000fffffffffffffff00000fffff"),
                (x"ffc0000000fffffffffffffe000000fffff"),
                (x"fffe000000fffffffffffffe000000fffff"),
                (x"fffe000000f8000003fffffe00001ffffff"),
                (x"fffe00000000000003ff000000001ffffff"),
                (x"fffe00000000000003ff000000001ffffff"),
                (x"fffe000000000000001f00000003fffffff"),
                (x"fffe000000000000000000000003fffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff800000000f800000000ffffffffff"),
                (x"ffffffffe000000f80000001fffffffffff"),
                (x"ffffffffe000000f80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 56_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffe000000fffffffffffffffffffffffff"),
                (x"fffe000000fffffffffffffffffffffffff"),
                (x"fffe00000007ffffffe000000ffffffffff"),
                (x"fffe000000003fffffe000000ffffffffff"),
                (x"fffffffc00003fffffe000000ffffffffff"),
                (x"fffffffc00003fffffe000000ffffffffff"),
                (x"fffffffc00003ffffc0000000ffffffffff"),
                (x"fffffffc00003fff800000000ffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffe00000000000fffffffffffffff"),
                (x"fffffffc000000000000fffffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff8000003ff0000007fffffffffffff"),
                (x"fffe00000007ffff80000001fffffffffff"),
                (x"fffe00000007ffff80000001fffffffffff"),
                (x"fffe00000007ffff80000001fffffffffff"),
                (x"fffe000000fffffffc0000000ffffffffff"),
                (x"fffe000000fffffffc0000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 57_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc0007fffffffffffff00000fffff"),
                (x"fffffffc0000000ffffffffe000000fffff"),
                (x"fffffffc0000000003fffffe000000fffff"),
                (x"fffffffc0000000003fffffe00001ffffff"),
                (x"ffffffffe0000000001ffffe00001ffffff"),
                (x"ffffffffe0000000001ffffe00001ffffff"),
                (x"fffffffffff800000000f8000003fffffff"),
                (x"fffffffffff80000000000000003fffffff"),
                (x"ffffffffffffc000000000000003fffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"ffffffffffffffff800000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffff800000000ffffffffff"),
                (x"ffffffffffffffff800000000ffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffff00000ffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 58_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffff000000001ffffff"),
                (x"fffe00000007fff00000000000001ffffff"),
                (x"ffc00000000000000000000000001ffffff"),
                (x"ffc00000000000000000000000001ffffff"),
                (x"ffc00000000000000000000000001ffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 59_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000f800007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"fffffffffff800007ffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 60_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffc00003fffffffffffffffffffffffffff"),
                (x"ffc00003fffffffffffffffffffffffffff"),
                (x"f8000003fffffffffffffffffffffffffff"),
                (x"f80000001ffffffffffffffffffffffffff"),
                (x"ffc0000000fffffffffffffffffffffffff"),
                (x"ffc0000000fffffffffffffffffffffffff"),
                (x"fffe00000007fffffffffffffffffffffff"),
                (x"fffe000000003ffffffffffffffffffffff"),
                (x"fffe000000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffff80000001fffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 61_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 62_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc0007fffffc0000000ffffffffff"),
                (x"fffffffc0007fffffc0000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 63_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"ffc0000000000000000000000000000001f"),
                (x"ffc0000000000000000000000000000001f"),
                (x"f800000000000000000000000000000001f"),
                (x"f800000000000000000000000000000001f"),
                (x"ffc000000000000003fffffffffffffffff"),

                -- 64_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 65_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffe000000003e000000ffffffffff"),
                (x"ffffffffe00000007fe000000ffffffffff"),
                (x"fffffffc0000000fffe000000ffffffffff"),
                (x"fffffffc000000007c000000007ffffffff"),
                (x"fffffffc000000007c000000007ffffffff"),
                (x"fffffffc000000007c000000007ffffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"ffffffffff000000000000000003fffffff"),
                (x"fffffffffff80000000000000003fffffff"),
                (x"ffffffffffffc000000000000003fffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 66_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe0000000001f0000007ffffffff"),
                (x"ffffffffe0003fffffff0000007ffffffff"),
                (x"ffffffffe0003fffffff0000007ffffffff"),
                (x"ffffffffe0003fffffff0000007ffffffff"),
                (x"ffffffffe0003fffffff0000007ffffffff"),
                (x"ffffffffe0003ff000000000007ffffffff"),
                (x"ffffffffe0003ff000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffff0000007ffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 67_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000ffffffffffffffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 68_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffff80000000007ffffffff"),
                (x"ffffffffffffc00000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffe0000000001f00000ffffffffff"),
                (x"ffffffffe00000007fff0000007ffffffff"),
                (x"fffffffc0000000fffe00000007ffffffff"),
                (x"fffffffc0000000fffe00000007ffffffff"),
                (x"fffffffc000000007fe000000ffffffffff"),
                (x"fffffffc000000007fe000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 69_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffe000000003ff0000007ffffffff"),
                (x"ffffffffe000000003ff0000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffe0000000001f0000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 70_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffffffff0000000000ffffffffff"),
                (x"fffffffffffffff0000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffc000001f0001fffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 71_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff80000000007fffffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"fffffffc0000000fffe000000ffffffffff"),
                (x"fffffffc0000000fffe000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffffffffffffff00000ffffffffff"),
                (x"ffffffffff00000ffc0000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 72_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff8000003fffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 73_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff003fffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 74_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffc0007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"ffffffffffffffff800007fffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc000001fffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),

                -- 75_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffffffffffffffffffff"),
                (x"ffffff8000fffffffc0007fffffffffffff"),
                (x"ffffff8000ffffff80000001fffffffffff"),
                (x"ffffff8000ffc00000000001fffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff8000000000001ffffffffffffffff"),
                (x"ffffff80000000000000fffffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff8000ffc00000000001fffffffffff"),
                (x"ffffff8000fffff0000000000ffffffffff"),
                (x"ffffff8000fffff0000000000ffffffffff"),
                (x"ffffff8000ffffff80000000007ffffffff"),
                (x"ffffff8000ffffffffe00000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007fffffffff800007ffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 76_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 77_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffe00000000000fffe0003fffffff"),
                (x"ffffffffe00000000000f80000001ffffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc0000000003ff000000000000000fffff"),
                (x"ffc0000000003ff000000001f00000fffff"),
                (x"ffc0000000003ff000000001f00000fffff"),
                (x"ffc0000000fffff0000007fff00000fffff"),
                (x"ffc0000000fffff0000007fff00000fffff"),
                (x"ffc0000000fffff0000007fff00000fffff"),
                (x"fffe000000fffff0000007fff00000fffff"),
                (x"fffe000000fffff0000007fff00000fffff"),
                (x"fffe000000fffff00000fffff00000fffff"),
                (x"fffe000000fffff00000fffff00000fffff"),
                (x"fffe000000fffff00000fffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffe000000fffffffffffffff00000fffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 78_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff800007fff00000fffffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff8000000000000007fffffffffffff"),
                (x"ffffff800000000000000001fffffffffff"),
                (x"ffffff800000000f80000001fffffffffff"),
                (x"ffffff8000003ffffc000001fffffffffff"),
                (x"ffffff8000003ffffc000001fffffffffff"),
                (x"ffffff8000003fffffe000000ffffffffff"),
                (x"ffffff8000003fffffe000000ffffffffff"),
                (x"ffffff8000003fffffe000000ffffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffff00000ffffffffff"),
                (x"ffffffffe0003ffffffffffffffffffffff"),
                (x"ffffffffe0003ffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 79_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffe00000007fe000000003fffffff"),
                (x"fffffffc000000007fff00000003fffffff"),
                (x"fffffffc0000000ffffff8000003fffffff"),
                (x"fffffffc00003ffffffff8000003fffffff"),
                (x"fffffffc00003ffffffff8000003fffffff"),
                (x"fffffffc0000000ffffff8000003fffffff"),
                (x"fffffffc0000000ffffff8000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 80_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffc00000000000007fffffffffffff"),
                (x"fffffffc0000000000000001fffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00003fff800000000ffffffffff"),
                (x"fffffffc00003ffffc000000007ffffffff"),
                (x"fffffffc00003fffffff00000003fffffff"),
                (x"fffffffc00003fffffff00000003fffffff"),
                (x"fffffffc00003fff800000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"fffffffc00003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff8000003ffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),

                -- 81_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000ffc000000007ffffffff"),
                (x"ffffffffe000000ffc000000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe000000fffff0000007ffffffff"),
                (x"ffffffffe00000007fe00000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffff00000000000000007ffffffff"),
                (x"ffffffffffffc00003e000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000ffffffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"ffffffffffffffffffe000000003fffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 82_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc00003ff0000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"ffffffffe000000ffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 83_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff000000000000000ffffffffff"),
                (x"ffffffffff0000007fff0001fffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"fffffffffff8000000000000007ffffffff"),
                (x"ffffffffffffc00000000000007ffffffff"),
                (x"ffffffffffffffffffe00000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffffffffffffff0000007ffffffff"),
                (x"ffffffffe000000ffc000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"ffffffffff00000000000001fffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 84_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 85_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000ffffffffff00000ffffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff8000003fffffe00000007ffffffff"),
                (x"ffffff800000000ffc000000007ffffffff"),
                (x"ffffff800000000ffc000000007ffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffe000000000000001fffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 86_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"ffffff8000003fffffff0000007ffffffff"),
                (x"ffffff8000003fffffff0000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc00003fffffe00000007ffffffff"),
                (x"fffffffc0000000ffc0000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffe0000000000007fffffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffff0000000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 87_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffc000001ffffffffffffffffffffffffff"),
                (x"ffc0000000ffffffffffffffff8000003ff"),
                (x"ffc0000000fffffffffffffff00000003ff"),
                (x"ffc0000000fffffffffffffff00000003ff"),
                (x"fffe00000007fffffffffffff00000fffff"),
                (x"fffe00000007fffffffffffff00000fffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff800007fffffffffffe00001ffffff"),
                (x"ffffff8000000000001ff80000001ffffff"),
                (x"ffffff8000000000001f000000001ffffff"),
                (x"fffffffc00000000000000000003fffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffffffe00000007c0000000ffffffffff"),
                (x"ffffffffffffffffffe00001fffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 88_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff800007fffffffffffffffffffffff"),
                (x"ffffff800000000ffffff800007ffffffff"),
                (x"ffffff800000000fffe00000007ffffffff"),
                (x"ffffff80000000007c000000007ffffffff"),
                (x"ffffff80000000007c000000007ffffffff"),
                (x"ffffffffe000000000000000007ffffffff"),
                (x"fffffffffff80000000000000ffffffffff"),
                (x"ffffffffff000000000007fffffffffffff"),
                (x"ffffffffe0000000000000000ffffffffff"),
                (x"fffffffc00000000000000000ffffffffff"),
                (x"ffffff80000000007fe00000007ffffffff"),
                (x"ffffff80000000007fe00000007ffffffff"),
                (x"ffffff8000003fffffe00000007ffffffff"),
                (x"ffffff800007ffffffe00000007ffffffff"),
                (x"ffffff800007ffffffff0000007ffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 89_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffff0001ffffff"),
                (x"fffffffc0000000ffffffffe00001ffffff"),
                (x"fffffffc0000000003fff80000001ffffff"),
                (x"fffffffc00000000001f000000001ffffff"),
                (x"fffffffc00000000001f000000001ffffff"),
                (x"ffffffffe0000000000000000003fffffff"),
                (x"ffffffffffffc00000000000007ffffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"ffffffffffffffff80000000007ffffffff"),
                (x"fffffffffffffffffc000000007ffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"fffffffffffffffffc0000000ffffffffff"),
                (x"ffffffffffffffff800000000ffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"fffffffffff800000000fffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff800007ffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 90_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff8000000000000000000ffffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffc0000000000000000007ffffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff800000000000000000007ffffffff"),
                (x"ffffff800000000ffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 91_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"ffffff800000000003fffffffffffffffff"),
                (x"ffffff800000000003fffffffffffffffff"),
                (x"ffffff80000000007ffffffffffffffffff"),
                (x"ffffff80000000007ffffffffffffffffff"),
                (x"ffffffffe00000007ffffffffffffffffff"),
                (x"ffffffffe000000003fffffffffffffffff"),
                (x"ffffffffff00000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000003fffffffffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"fffffffffff8000000000001fffffffffff"),
                (x"ffffffffffffc00000000001fffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 92_character
                (x"ffffffffffffc00003fffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 93_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"fffffffc0000000003fffffffffffffffff"),
                (x"fffffffc00000000001ffffffffffffffff"),
                (x"fffffffc00000000001ffffffffffffffff"),
                (x"ffffffffe0000000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff00000fffffffffffffff"),
                (x"fffffffffffffff0000007fffffffffffff"),
                (x"fffffffffffffff000000001fffffffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"fffffffffffffff000000000007ffffffff"),
                (x"ffffffffffffffff80000000007ffffffff"),
                (x"ffffffffffffffff80000000007ffffffff"),
                (x"ffffffffffffc00000000000007ffffffff"),
                (x"ffffffffffffc000000000000ffffffffff"),
                (x"ffffffffffffc000000007fffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc0000000fffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"ffffffffffffc000001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffffffff0001ffffffffffffffff"),
                (x"fffffffffff80000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"ffffffffff000000001ffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 94_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffffffffe000000003fffffff0001ffffff"),
                (x"ffffff8000000000001ffffe00001ffffff"),
                (x"fffe0000000000000000fffe00001ffffff"),
                (x"ffc00000000000000000000000001ffffff"),
                (x"ffc00000000000000000000000001ffffff"),
                (x"ffc0000000ffc0000000000000001ffffff"),
                (x"ffc0000000fffff00000000000001ffffff"),
                (x"ffc000001fffffff800000000003fffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),

                -- 95_character
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"ffc00003fffffffffffffffffffffffffff"),
                (x"ffc000000000000000000000007ffffffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc000000000000000000000000000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc00003fffffffffffffffff00000fffff"),
                (x"ffc000001ffffffffffffffff00000fffff"),
                (x"ffc000001fffffffffffffffff8000fffff"),
                (x"ffc000001fffffffffffffffff8000003ff"),
                (x"ffc000001fffffffffffffffff8000003ff"),
                (x"ffc000001fffffffffffffffff8000003ff"),
                (x"ffc000001fffffffffffffffff8000003ff"),
                (x"ffc000001fffffffffffffffff8000003ff"),
                (x"ffc000001fffffffffffffffff80000001f"),
                (x"ffc000001fffffffffffffffff80000001f"),
                (x"ffc000001ffffffffffffffffffc000001f"),
                (x"ffc000001ffffffffffffffffffc000001f"),
                (x"ffc000001ffffffffffffffffffc000001f"),
                (x"ffc000001ffffffffffffffffffc000001f"),
                (x"ffc000001ffffffffffffffffffc000001f"),
                (x"ffc0000000000000000000000000000001f"),
                (x"ffc0000000000000000000000000000001f"),
                (x"ffc000000000000000000000000000003ff"),
                (x"ffc000000000000000000000000000003ff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff"),
                (x"fffffffffffffffffffffffffffffffffff")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 3551 := 0;
    signal out_color_reg : std_logic_vector(139 downto 0) := (others => '0');
begin
    process(in_sprite_id, in_sprite_row, in_sprite_col, in_sprite_state, in_sprite_direction)
    begin
        real_row <= 0;
        case in_sprite_id is
            when 0 => real_row <= in_sprite_row;
            when 1 => real_row <= 37 + in_sprite_row;
            when 2 => real_row <= 74 + in_sprite_row;
            when 3 => real_row <= 111 + in_sprite_row;
            when 4 => real_row <= 148 + in_sprite_row;
            when 5 => real_row <= 185 + in_sprite_row;
            when 6 => real_row <= 222 + in_sprite_row;
            when 7 => real_row <= 259 + in_sprite_row;
            when 8 => real_row <= 296 + in_sprite_row;
            when 9 => real_row <= 333 + in_sprite_row;
            when 10 => real_row <= 370 + in_sprite_row;
            when 11 => real_row <= 407 + in_sprite_row;
            when 12 => real_row <= 444 + in_sprite_row;
            when 13 => real_row <= 481 + in_sprite_row;
            when 14 => real_row <= 518 + in_sprite_row;
            when 15 => real_row <= 555 + in_sprite_row;
            when 16 => real_row <= 592 + in_sprite_row;
            when 17 => real_row <= 629 + in_sprite_row;
            when 18 => real_row <= 666 + in_sprite_row;
            when 19 => real_row <= 703 + in_sprite_row;
            when 20 => real_row <= 740 + in_sprite_row;
            when 21 => real_row <= 777 + in_sprite_row;
            when 22 => real_row <= 814 + in_sprite_row;
            when 23 => real_row <= 851 + in_sprite_row;
            when 24 => real_row <= 888 + in_sprite_row;
            when 25 => real_row <= 925 + in_sprite_row;
            when 26 => real_row <= 962 + in_sprite_row;
            when 27 => real_row <= 999 + in_sprite_row;
            when 28 => real_row <= 1036 + in_sprite_row;
            when 29 => real_row <= 1073 + in_sprite_row;
            when 30 => real_row <= 1110 + in_sprite_row;
            when 31 => real_row <= 1147 + in_sprite_row;
            when 32 => real_row <= 1184 + in_sprite_row;
            when 33 => real_row <= 1221 + in_sprite_row;
            when 34 => real_row <= 1258 + in_sprite_row;
            when 35 => real_row <= 1295 + in_sprite_row;
            when 36 => real_row <= 1332 + in_sprite_row;
            when 37 => real_row <= 1369 + in_sprite_row;
            when 38 => real_row <= 1406 + in_sprite_row;
            when 39 => real_row <= 1443 + in_sprite_row;
            when 40 => real_row <= 1480 + in_sprite_row;
            when 41 => real_row <= 1517 + in_sprite_row;
            when 42 => real_row <= 1554 + in_sprite_row;
            when 43 => real_row <= 1591 + in_sprite_row;
            when 44 => real_row <= 1628 + in_sprite_row;
            when 45 => real_row <= 1665 + in_sprite_row;
            when 46 => real_row <= 1702 + in_sprite_row;
            when 47 => real_row <= 1739 + in_sprite_row;
            when 48 => real_row <= 1776 + in_sprite_row;
            when 49 => real_row <= 1813 + in_sprite_row;
            when 50 => real_row <= 1850 + in_sprite_row;
            when 51 => real_row <= 1887 + in_sprite_row;
            when 52 => real_row <= 1924 + in_sprite_row;
            when 53 => real_row <= 1961 + in_sprite_row;
            when 54 => real_row <= 1998 + in_sprite_row;
            when 55 => real_row <= 2035 + in_sprite_row;
            when 56 => real_row <= 2072 + in_sprite_row;
            when 57 => real_row <= 2109 + in_sprite_row;
            when 58 => real_row <= 2146 + in_sprite_row;
            when 59 => real_row <= 2183 + in_sprite_row;
            when 60 => real_row <= 2220 + in_sprite_row;
            when 61 => real_row <= 2257 + in_sprite_row;
            when 62 => real_row <= 2294 + in_sprite_row;
            when 63 => real_row <= 2331 + in_sprite_row;
            when 64 => real_row <= 2368 + in_sprite_row;
            when 65 => real_row <= 2405 + in_sprite_row;
            when 66 => real_row <= 2442 + in_sprite_row;
            when 67 => real_row <= 2479 + in_sprite_row;
            when 68 => real_row <= 2516 + in_sprite_row;
            when 69 => real_row <= 2553 + in_sprite_row;
            when 70 => real_row <= 2590 + in_sprite_row;
            when 71 => real_row <= 2627 + in_sprite_row;
            when 72 => real_row <= 2664 + in_sprite_row;
            when 73 => real_row <= 2701 + in_sprite_row;
            when 74 => real_row <= 2738 + in_sprite_row;
            when 75 => real_row <= 2775 + in_sprite_row;
            when 76 => real_row <= 2812 + in_sprite_row;
            when 77 => real_row <= 2849 + in_sprite_row;
            when 78 => real_row <= 2886 + in_sprite_row;
            when 79 => real_row <= 2923 + in_sprite_row;
            when 80 => real_row <= 2960 + in_sprite_row;
            when 81 => real_row <= 2997 + in_sprite_row;
            when 82 => real_row <= 3034 + in_sprite_row;
            when 83 => real_row <= 3071 + in_sprite_row;
            when 84 => real_row <= 3108 + in_sprite_row;
            when 85 => real_row <= 3145 + in_sprite_row;
            when 86 => real_row <= 3182 + in_sprite_row;
            when 87 => real_row <= 3219 + in_sprite_row;
            when 88 => real_row <= 3256 + in_sprite_row;
            when 89 => real_row <= 3293 + in_sprite_row;
            when 90 => real_row <= 3330 + in_sprite_row;
            when 91 => real_row <= 3367 + in_sprite_row;
            when 92 => real_row <= 3404 + in_sprite_row;
            when 93 => real_row <= 3441 + in_sprite_row;
            when 94 => real_row <= 3478 + in_sprite_row;
            when 95 => real_row <= 3515 + in_sprite_row;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= rom(real_row);
        end if;
    end process;
    out_color <= out_color_reg(((in_sprite_col + 1) * 5) - 1 downto (in_sprite_col * 5));
end behavioral;
