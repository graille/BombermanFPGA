library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.PROJECT_PARAMS_PKG.all;
use work.PROJECT_TYPES_PKG.all;
use work.PROJECT_DIRECTION_PKG.all;

entity sprite_rom is
    port (
        clk : in std_logic;

        in_sprite_id : in block_category_type;
        in_sprite_state : in state_type;
        in_sprite_direction : in direction_type;
        in_sprite_row : in integer range 0 to 51;
        in_sprite_col : in integer range 0 to 49;

        out_color : out std_logic_vector(4 downto 0) := (others => '0')
    );
end sprite_rom;

architecture behavioural of sprite_rom is
    subtype word_t is std_logic_vector(49 downto 0);
    type memory_t is array(2051 downto 0) of word_t;

    function init_mem 
        return memory_t is
        begin
            return (
                -- 1_unbreakable
                ("1110111101111010111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110010000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010000100000110001100011011110111101111"),
                ("1110111101111010111101111011110010000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010000100000110001100011011110111101111"),
                ("1110111101111010111101111011110010000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010000100000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110000100001000010000100001000010010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000001000010000100001000010000100001000110001100011011110111101111"),
                ("1110111101111010111101111011110010000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010000100000110001100011011110111101111"),
                ("1110111101111010111101111011110010000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010000100000110001100011011110111101111"),
                ("1110111101111010111101111011110010000100001000000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001000010000100000110001100011011110111101111"),
                ("1110111101111010111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011011110111101111"),
                ("1110111101111010111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011011110111101111"),
                ("1110111101111010111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011011110111101111"),
                ("1110111101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("1110111101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("1110111101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("1110111101111011111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111"),
                ("1110111101111011110111101111011111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110"),
                ("1110111101111011110111101111011111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110"),
                ("1110111101111011110111101111011111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110"),
                ("1110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111101111011110"),
                ("1110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111101111011110"),
                ("1110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111101111011110"),
                ("1110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100"),
                ("1110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100"),
                ("1110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100"),

                -- 2_unbreakable
                ("1110011100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("1110011100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("1110011100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("1110011100111000111101111011110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000110001100011111011110111101"),
                ("1110011100111000111101111011110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000110001100011111011110111101"),
                ("1110011100111000111101111011110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000110001100011111011110111101"),
                ("1110011100111001111011110111100001100011000110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100001100011000110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100001100011000110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001101111011110111100100001000010000011000110001100011000110001101111011110111100100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001101111011110111100100001000010000011000110001100011000110001101111011110111100100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001101111011110111100100001000010000011000110001100011000110001101111011110111100100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100100001000010000100001000010000011000110001100011000110001100100001000010000100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001101111011110111100100001000010000011000110001100011000110001101111011110111100100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001101111011110111100100001000010000011000110001100011000110001101111011110111100100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001101111011110111100100001000010000011000110001100011000110001101111011110111100100001000010001111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001101111011110111100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111111011110111101"),
                ("1110011100111001111011110111100111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111111011110111101"),
                ("1110011100111001111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110011110111101111111011110111101"),
                ("1110011100111001111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110011110111101111111011110111101"),
                ("1110011100111001111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110011110111101111111011110111101"),
                ("1110011100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("1110011100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("1110011100111001110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111101"),
                ("1110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111011110111101"),
                ("1110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111011110111101"),
                ("1110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111011110111101"),

                -- 3_breakable
                ("0011000110001100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100011000111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011000110001100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100011000111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011000110001100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100011000111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100011000111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100011000111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000110001100011000111001110011100011000110001100011000110001100011000110001100011000110001100011"),
                ("0011100111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100110001100011000111001110011100111001110011100111001110011100111001110011100111001110011100111"),
                ("0011100111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100110001100011000111001110011100111001110011100111001110011100111001110011100111001110011100111"),
                ("0011100111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100110001100011000111001110011100111001110011100111001110011100111001110011100111001110011100111"),
                ("0011100111001110010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100110001100011000111001110011100111001110011100111001110011100111001110011100111001110011100111"),
                ("0011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("0011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("0011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("0010100101001010010100101001010010100101001010011000110001100010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000110000110001100011001010010100101"),
                ("0010100101001010010100101001010010100101001010011000110001100010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000110000110001100011001010010100101"),
                ("0010100101001010010100101001010010100101001010011000110001100010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001100011000110000110001100011001010010100101"),
                ("0010100101001010010100101001010010100101001010011000110001100010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111000110001100011001010010100101"),
                ("0010100101001010010100101001010010100101001010011000110001100010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111000110001100011001010010100101"),
                ("0010100101001010010100101001010010100101001010011000110001100010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111000110001100011001010010100101"),
                ("0001100011000110001100011000110001100011000110011100111001110010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111000110001100011000110001100011"),
                ("0001100011000110001100011000110001100011000110011100111001110010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111000110001100011000110001100011"),
                ("0001100011000110001100011000110001100011000110011100111001110010100101001010010100100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001110011100111000110001100011000110001100011"),
                ("0001100011000110001100011000110001100011000110011000110001100010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001110011100111000110001100011000110001100011"),
                ("0001100011000110001100011000110001100011000110011000110001100010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001110011100111000110001100011000110001100011"),
                ("0001100011000110001100011000110001100011000110011000110001100010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001110011100111000110001100011000110001100011"),
                ("0011100111001110011000110001100011000110001100011000110001100011000110001100011000111001110011100110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001110011100111001110011100111001110011100111"),
                ("0011100111001110011000110001100011000110001100011000110001100011000110001100011000111001110011100110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001110011100111001110011100111001110011100111"),
                ("0011100111001110011000110001100011000110001100011000110001100011000110001100011000111001110011100110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001110011100111001110011100111001110011100111"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001000010000100001000010000100001000010000100"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100111001110011100011000110001100011000110001100011000110001100011000110001100011000110001100110001100011000110001010010100101001010010100101001010010100101"),
                ("0011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001110011100111001110011100111001110011100111"),
                ("0011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001110011100111001110011100111001110011100111"),
                ("0011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110001100011000110001110011100111001110011100111001110011100111"),
                ("0011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("0011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),
                ("0011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110001100011000110"),

                -- 4_bomb_0
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000100001000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000100001000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000100001000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000100111001110011010000100001000111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000100111001110011010000100001000111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000100111001110011010000100001000111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001110011100111001110011100111001110011100111001110011100111001110011100111111111111111000000000000000111111111111111000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001110011100111001110011100111001110011100111001110011100111001110011100111111111111111000000000000000111111111111111000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001110011100111001110011100111001110011100111001110011100111001110011100111111111111111000000000000000111111111111111000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110000000000000000011000110001100011000110001100000100001000010011000110001101110011100111001110011100000010000100001000000000000000111111111111111000000000000000000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110000000000000000011000110001100011000110001100000100001000010011000110001101110011100111001110011100000010000100001000000000000000111111111111111000000000000000000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111110000000000000000011000110001101000110001100011000110001100011000110001100010011000110001100011000110111001110011100000010000100001000000000000000000000000000000111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000000011000110001101000110001100011000110001100011000110001100010011000110001100011000110111001110011100000010000100001000000000000000000000000000000111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000000011000110001101000110001100011000110001100011000110001100010011000110001100011000110111001110011100000010000100001000000000000000000000000000000111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001000110001100010000100001000010000100001000010101101011010111000110001100010011000110111001110011100111111111111111111111111111111111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001000110001100010000100001000010000100001000010101101011010111000110001100010011000110111001110011100111111111111111111111111111111111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001000110001100010000100001000010000100001000010101101011010111000110001100010011000110111001110011100111111111111111111111111111111111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111110000000000000000011000110001101000110001100010000100001000010000100001000010101101011010111000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100010000100001000010000100001000010101101011010111000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100010000100001000010000100001000010101101011010111000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100010101101011010110101101011010110101101011010111000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100010101101011010110101101011010110101101011010111000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100010101101011010110101101011010110101101011010111000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100011000110001100011000110001100011000110001100011000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100011000110001100011000110001100011000110001100011000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001101000110001100011000110001100011000110001100011000110001100011000110001100010011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001100011000110001101000110001100011000110001100011000110001100010011000110001100011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001100011000110001101000110001100011000110001100011000110001100010011000110001100011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000000011000110001100011000110001101000110001100011000110001100011000110001100010011000110001100011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000001110011100111000011000110001100011000110001100011000110001100011000110001100011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000001110011100111000011000110001100011000110001100011000110001100011000110001100011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000001110011100111000011000110001100011000110001100011000110001100011000110001100011000110001100011000110111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000001110011100111001110011100111000011000110001100011000110001100011000110001101110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000001110011100111001110011100111000011000110001100011000110001100011000110001101110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111110000000000000001110011100111001110011100111000011000110001100011000110001100011000110001101110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000"),
                ("1111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111"),
                ("1111111111111111111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000000000000000000111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000000000000000000111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001110011100111001110011100111001110011100111001110011100111001110011100111001110011100000000000000000000000000000000111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 5_explosion_0
                ("1111111111111111111111111111110110001100110011100111001101101011011010010010100101001010010100111000101101011010011010010100101001010010100110011100111001110110101101001111001110011100111001110011100111001110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001101101011011010010010100101001010010100111000101101011010011010010100101001010010100110011100111001110110101101001111001110011100111001110011100111001110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100110011110101101011000110001100011000100111001110110110101101001001010010100111010110101101010011100111011011001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001101101011010011100111001110110101101011010011010010100101001010011100011000110001100010011100111011010011100111001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001101101011010011100111001110110101101011010011010010100101001010011100011000110001100010011100111011010011100111001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111011001100111001110011100111001110011100110011101101011010110101101011010011110101101001001010010100101001010010100101001010011101010110101101011010110101101100111001110011100111001110011100111001110011111111111111111111111111"),
                ("1111011110111101111011110011001100111001110011100111001100111001110110101101011010110101101011011010010010100111010110101101001001010011101011010110101101010011100111001111001110011100111001110011100111001110011100111001110010110001100011001100111001"),
                ("1111011110111101111011110011001100111001110011100111001100111001110110101101011010110101101011011010010010100111010110101101001001010011101011010110101101010011100111001111001110011100111001110011100111001110011100111001110010110001100011001100111001"),
                ("0111001110011100110001100110011100111001110011100111001100111001110110101101011010110101101011011010010010100111000010010100101001010011100011010110101001110110101101100111001110011011010011100111001110011110011100111001110011100111001100110110001100"),
                ("1110111101011001100111001100111100111001110011100111001100111001111001100111001111001100111001111000110101101011010010010100101001010010100110011100111011010110101101001111001110011011010110101101100111001110011100111001110011001110011100110110001100"),
                ("1110111101011001100111001100111100111001110011100111001100111001111001100111001111001100111001111000110101101011010010010100101001010010100110011100111011010110101101001111001110011011010110101101100111001110011100111001110011001110011100110110001100"),
                ("1100111001110011100111001100111011010110110011001110011100111001111001110011100111001100111001111000110101101010011110101101001001010010100111010110101101010011100111001110011100111100110011100111001110011110011100111001100111011010110110011100111001"),
                ("1100111001110011100111001100111011010110110011001110011100111001111001110011100111001100111001111000110101101010011110101101001001010010100111010110101101010011100111001110011100111100110011100111001110011110011100111001100111011010110110011100111001"),
                ("1100111001110011100111001110011100111001100111011010110101101011010110100111001111001100111001111000110001100011010110001100001001010010100111000110000100111010110101011010110101101001110011100111011010110100111001110011110011100111001110011001110011"),
                ("1100111001110011100111001110011011010110101101011010110101101011010011100111001110011110101101001001010010100101001010010100101001010010100101001010010100111010110101011010011100111011010110101101011010110101101011010110100111001110011100111011010110"),
                ("1100111001110011100111001110011011010110101101011010110101101011010011100111001110011110101101001001010010100101001010010100101001010010100101001010010100111010110101011010011100111011010110101101011010110101101011010110100111001110011100111011010110"),
                ("1101011010110101001110011100111011010110101101011010110101101011011010110001100010011110101101011010110001100001001010010100101001010010100101001010010100101001010011100010011100111011010110101101011010110101101011010110101101011010110101101011010110"),
                ("0100101001110001001110011101101011010110101101011010110100111001111010101101011010011010010100101001110101101011010010010100111000110000100101001010010100101001010011101010011100111011010110101101011010110101101001110011100111001110011101101011010110"),
                ("0100101001110001001110011101101011010110101101011010110100111001111010101101011010011010010100101001110101101011010010010100111000110000100101001010010100101001010011101010011100111011010110101101011010110101101001110011100111001110011101101011010110"),
                ("0100101001110101001110011101101001110011101101011010110100111001111010101101011010110110101101001001110001100001000010010100101001010010100101001010010100111000110001001110011100111011010011100111011010110100111100011000110001100011000110100110001100"),
                ("0100101001110101001110011100111001110011100111011010110101101011011000110101101010110100111001111000010010100101000010000100001001010010100101001010010100111000110001001111010110101101011010110101011010110100111100011000010010100101001010011111011110"),
                ("0100101001110101001110011100111001110011100111011010110101101011011000110101101010110100111001111000010010100101000010000100001001010010100101001010010100111000110001001111010110101101011010110101011010110100111100011000010010100101001010011111011110"),
                ("0100101001110101011010110101101011010110100111001110011100111001111000110001100011010110101101011010010010100101000010010100101001010010100101001010010100111000110000100101000010000100111000110000100101001110101101011010010010100101001010011101011010"),
                ("0100101001010011001110011101101011010110100110100101001010010100111000110001100001001010010100111000010010100101001110001100001001010010100001001010011100001001010010100001000010000100101001010010100101001110101101011010010011100011000010011100011000"),
                ("0100101001010011001110011101101011010110100110100101001010010100111000110001100001001010010100111000010010100101001110001100001001010010100001001010011100001001010010100001000010000100101001010010100101001110101101011010010011100011000010011100011000"),
                ("1100011000110000100101001010000100001000100111100011000010010100101001010010100101001010010100101001110001100011000010010100101001010010100001001010010100111000110001101001001010010100101001010011101011010110100100101001110101100011000010010100101001"),
                ("1100011000110000100101001010000100001000100111100011000010010100101001010010100101001010010100101001110001100011000010010100101001010010100001001010010100111000110001101001001010010100101001010011101011010110100100101001110101100011000010010100101001"),
                ("0100101001010010100101001010000100101001010000100101001110001100001001010000100001001110101101001001110001100001001010000100001000010000100101001010010100110011100111001111010110101101010011100111001110011110101100011000100111101011010110100100101001"),
                ("0100101001010010100101001110001101011010010011101011010110001100001001010010100110011100111001101001110001100001001010000100001000010000100001001010010100001001010011101010011100111001110011100111011010110100111001110011100110100101001110000100101001"),
                ("0100101001010010100101001110001101011010010011101011010110001100001001010010100110011100111001101001110001100001001010000100001000010000100001001010010100001001010011101010011100111001110011100111011010110100111001110011100110100101001110000100101001"),
                ("1100011000010011101011010100111011010110101101001110011010010100101001010010100111010100111001101001010010100101001010010100101000010000100101001010010100101001010010100111000110001001111000110001001110011101101011010110100111001110011010011101011010"),
                ("0100101001010011101011010101101011010110101101001110011100111001110011110101101011010110101101011000010010100101001010010100101001010011100001001010011100001001010010100101001010011101010011100111011010110101101011010110110011100111001100111100011000"),
                ("0100101001010011101011010101101011010110101101001110011100111001110011110101101011010110101101011000010010100101001010010100101001010011100001001010011100001001010010100101001010011101010011100111011010110101101011010110110011100111001100111100011000"),
                ("1101011010100111011010110101101011010110101101011010110101101011010110101101011010110100111001101001010010100101001010010100101001010010100101001010010100101001010011101011010110101001110110101101011010110101101001110011110011011010110100111101011010"),
                ("1001110011101101011010110110011001110011101101011010110101101011010110101101011010110101101011011010110101101011000010010100101001010010100101001010011101010011100111011010110101101011010110101101011010110100111100111001100111001110011100111001110011"),
                ("1001110011101101011010110110011001110011101101011010110101101011010110101101011010110101101011011010110101101011000010010100101001010010100101001010011101010011100111011010110101101011010110101101011010110100111100111001100111001110011100111001110011"),
                ("1100111001110011011010110100111100111001100111011010110100111001110110101101011010011101101011010110100111001101001110001100011010110101101001001010011001110110101101011010110101101001110110101101001110011110011100111001101101001110011100111011010110"),
                ("0110001100110011100111001110011100111001110011100111001110011100111001110011100111001110011100110011110001100001001110001100010110101101011010011100111001111001110011001110110101101011010011100111100111001110011100111001110011001110011100111111011110"),
                ("0110001100110011100111001110011100111001110011100111001110011100111001110011100111001110011100110011110001100001001110001100010110101101011010011100111001111001110011001110110101101011010011100111100111001110011100111001110011001110011100111111011110"),
                ("0111001110111011100111001110011100111001110011100111001110011100111001110011100111001110011100110011010010100111000110101101010011100111001110011100111101011001110011100110011100111100111001110011100111001110011100111001110011100111001110010110001100"),
                ("0111001110111011100111001110011100111001110011100111001110011100111001110011100111001110011100110011010010100111000110101101010011100111001110011100111101011001110011100110011100111100111001110011100111001110011100111001110011100111001110010110001100"),
                ("1111011110111011100111001110011100111001110011100111001110011100110011100111001111001110011100111010010010100101001110001100011010110101101011010110101100010011100111011010110101101100111001110011100111001110011100111001110011100111001110011100111001"),
                ("1100111001110011100111001011001100111001110011100111001110011100111001101101011010110101101011010110110101101001001010010100101001010010100101001010011101010110101101011010011100111100111001110011100111001110011100111001110011100111001011000110001100"),
                ("1100111001110011100111001011001100111001110011100111001110011100111001101101011010110101101011010110110101101001001010010100101001010010100101001010011101010110101101011010011100111100111001110011100111001110011100111001110011100111001011000110001100"),
                ("1111111111111111111111111011001100111001110011100111001110011100111001101101011010110101101011010110100111001101001010010100101001010010100111010110101001110110101101011010110101101100111001110011100111001110011100111001110011111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001101101011010110101101011010110100111001110011110001100001000010000100010011100111001110011100111001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001101101011010110101101011010110100111001110011110001100001000010000100010011100111001110011100111001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110110011100111001110011100111001101101011010110101101011010110101101011010110100111001111000110000100111010110101001110011100111100111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111100110001100011001100111001110011100110011110011100110011110101101010011100111001110110110101101001000010000100101000010000100001001010011001111001110011100111001110011100111001110011100111001100111111111111111111111111111"),
                ("1111111111111111111111111111100110001100011001100111001110011100110011110011100110011110101101010011100111001110110110101101001000010000100101000010000100001001010011001111001110011100111001110011100111001110011100111001100111111111111111111111111111"),

                -- 5_explosion_1
                ("1100111001110011110111101111101100111001110011100111001110101101001001010010100111000010010100101001010010100101001010000100001000010000100001000010000100001001010011101011010110101101001001010011001110011101101011010110100111100111001111101111011110"),
                ("1100111001110011110111101111101100111001110011100111001110101101001001010010100111000010010100101001010010100101001010000100001000010000100001000010000100001001010011101011010110101101001001010011001110011101101011010110100111100111001111101111011110"),
                ("1100111001110010110001100111011100111001101101001110011010010100101001010010100101001110001100001001010000100001000010000100001000010000100001001010010100001001010010100111000110000100111010110101001110011100111011010110100111100111001011001100111001"),
                ("1001110011101101011010110100111001110011100111101011010010010100111000110001100011000110001100001001010000100001000010000100001000010000100001000010000100101000010000100111000110001101010011100111001110011100111011010110101101100111001110010110001100"),
                ("1001110011101101011010110100111001110011100111101011010010010100111000110001100011000110001100001001010000100001000010000100001000010000100001000010000100101000010000100111000110001101010011100111001110011100111011010110101101100111001110010110001100"),
                ("1011010110101101011010110101101011010110100111101011010110001100001001010010100101001010010100101001010000100001000010000100001000010000100001000010000100101001010010100111010110101101011000110001001110011100111011010110100111100111001110011100111001"),
                ("1011010110101101011010110101101001110011100111001110011110101101001001010010100101001010010100101000010000100001000010000100001000010000100001000010000100101001010011100011010110100100111000110001001110011100111011010110101101001110011100111001110011"),
                ("1011010110101101011010110101101001110011100111001110011110101101001001010010100101001010010100101000010000100001000010000100001000010000100001000010000100101001010011100011010110100100111000110001001110011100111011010110101101001110011100111001110011"),
                ("1011010110101101011010110101101101011010110101101011010010010100101001010010100111000010010100101001010010100101000010000100001000010000100001000010000100001001010011100011010110100100111000110001001110011100111011010110101101011010110101101001110011"),
                ("1001110011101101011010110101101001110011010010100101001010010100101001010010100101001110001100001001010000100001000010000100001000010000100001001010010100101001010010100101001010010100101001010010100101001100111011010110100111011010110100111001110011"),
                ("1001110011101101011010110101101001110011010010100101001010010100101001010010100101001110001100001001010000100001000010000100001000010000100001001010010100101001010010100101001010010100101001010010100101001100111011010110100111011010110100111001110011"),
                ("0100101001100111011010110100111011010110110100100101001010010100101001010010100101001110001100001001010000100001000010000100001000010000100111000110000100101001010010100101001010010100101001010010100101001110101101011010010011101011010110101001110011"),
                ("0100101001100111011010110100111011010110110100100101001010010100101001010010100101001110001100001001010000100001000010000100001000010000100111000110000100101001010010100101001010010100101001010010100101001110101101011010010011101011010110101001110011"),
                ("0100101001110101011010110110101101011010110000100101001010010100111000110001100011000110001100001001010000100001000010000100001000010000100111000110000100101001010011100011000110001100001001010010100101001010010100101001010010100101001110101001110011"),
                ("1100011000110001101011010110000100101001010010100101001110001100001001010010100101001010010100101000010000100001000010000100001000010000100101001010010100101001010010100101001010010100111000110000100101001010000100101001110001100011000010011100011000"),
                ("1100011000110001101011010110000100101001010010100101001110001100001001010010100101001010010100101000010000100001000010000100001000010000100101001010010100101001010010100101001010010100111000110000100101001010000100101001110001100011000010011100011000"),
                ("0100101001010010100101001010010100101001010010100101001010010100101001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110000100101001010000100101001010000100101001110000100101001"),
                ("0100101001010010100101001110001100011000010010100001000010010100101001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010000100001000010000100101001110000100001000"),
                ("0100101001010010100101001110001100011000010010100001000010010100101001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010000100001000010000100101001110000100001000"),
                ("0100101001010000100001000010010100101001010010100101001010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010001100001000010000100001000010000100001000010011101011010010010001100011"),
                ("0100101001010000100001000010000100001000010000100101001010010100101000010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001000"),
                ("0100101001010000100001000010000100001000010000100101001010010100101000010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100101001010010100101001010000100001000010000100001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100101001010010100101001010000100001000010000100001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100101001010010100001000010000100001000010010100101001110001100001001010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001"),
                ("0100001000110001100011000010010100001000010000100101001010010100101001110001100001001010000100001000010000100001000010000100001000010000100001000010000100101000010000100101001010010100101001010010100101001010000100001000010000100001000010000100001000"),
                ("0100001000110001100011000010010100001000010000100101001010010100101001110001100001001010000100001000010000100001000010000100001000010000100001000010000100101000010000100101001010010100101001010010100101001010000100001000010000100001000010000100001000"),
                ("0100101001010010100101001010010100101001010010100001000010000100001001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001010010100111000110001100011000010010100101001110000100101001010010100101001"),
                ("0100101001010010100101001010010100101001010010100101001010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100001000010000100101001110000100101001010011100011000110001100011000"),
                ("0100101001010010100101001010010100101001010010100101001010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100001000010000100101001110000100101001010011100011000110001100011000"),
                ("0100101001010010100101001110000100101001010010100101001010000100001000110001100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100111000110000100101000010000100101001110000100101001010010100101001010010100101001"),
                ("1101011010110000100101001010010100101001110001100011000010010100101001110001100011000110001100001001010000100001000010000100001000010000100001000010000100001000010000100101000010001100001001010010100101001010010100101001010010100101001010010100101001"),
                ("1101011010110000100101001010010100101001110001100011000010010100101001110001100011000110001100001001010000100001000010000100001000010000100001000010000100001000010000100101000010001100001001010010100101001010010100101001010010100101001010010100101001"),
                ("1101011010110100100101001010011100011000010010100101001110001100011000010010100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100101000010000100111000110000100101001010010100101001010011100011000100110100101001"),
                ("0100101001010011100011000010011101011010110000100101001010010100101001010010100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010010100101001010010100101001100111100011000"),
                ("0100101001010011100011000010011101011010110000100101001010010100101001010010100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010010100101001010010100101001100111100011000"),
                ("1101011010110101001110011010011100011000100111100011000010010100101001010010100111000110001100001001010010100101001010000100001000010000100001000010000100001001010010100101000010000100111000110001100011000010011100011000110101001110011101101001110011"),
                ("1101011010110101001110011010011100011000100111100011000010010100101001010010100111000110001100001001010010100101001010000100001000010000100001000010000100001001010010100101000010000100111000110001100011000010011100011000110101001110011101101001110011"),
                ("1001110011100111101011010010011100011000101101101011010010010100101001110001100001001010010100111000010010100101001010000100001000010000100001000010000100101001010010100001001010011100011000110001001110011100111101011010100111001110011100111011010110"),
                ("1011010110100111001110011100111001110011101101001110011010010100101001110101101001001010010100111000010010100101000010000100001000010000100001000010000100101000010000100001001010010100111000110001001110011101101011010110101101011010110101101011010110"),
                ("1011010110100111001110011100111001110011101101001110011010010100101001110101101001001010010100111000010010100101000010000100001000010000100001000010000100101000010000100001001010010100111000110001001110011101101011010110101101011010110101101011010110"),
                ("1001110011110011011010110101101011010110101101001110011110001100011000100111001110110110001100001001010010100111000010010100101000010000100001000010000100001001010011100011000110001101010011100111001110011101101011010110101101011010110100111001110011"),
                ("1100111001110011011010110100111011010110101101011010110110101101010011100111001110011110101101001001010010100111000010010100101000010000100001001010010100101001010010100001001010011100011000110001001110011101101001110011110011100111001110011100111001"),
                ("1100111001110011011010110100111011010110101101011010110110101101010011100111001110011110101101001001010010100111000010010100101000010000100001001010010100101001010010100001001010011100011000110001001110011101101001110011110011100111001110011100111001"),
                ("1100111001110011100111001110011001110011101101001110011100111001110110110101101001001110001100001001010010100101001010000100001000010000100001001010010100001000010000100001001010011100001001010011101011010101101100111001110011100111001110010110001100"),
                ("1100111001110011100111001110011100111001101101011010110101101011011000010010100101001110001100001001010000100001000010000100001000010000100001000010000100001000010000100001001010011100001001010011101011010101101100111001110011100111001111010111001110"),
                ("1100111001110011100111001110011100111001101101011010110101101011011000010010100101001110001100001001010000100001000010000100001000010000100001000010000100001000010000100001001010011100001001010011101011010101101100111001110011100111001111010111001110"),

                -- 5_explosion_2
                ("1111111111110010110001100110011100111001101101001110011110001100001001010000100001000010000100001000010000100001000010000100011011110111101101000010000100001000010000100111000110001101011000110001101011010101100110001100111100110001100111101111011110"),
                ("1111111111110010110001100110011100111001101101001110011110001100001001010000100001000010000100001000010000100001000010000100011011110111101101000010000100001000010000100111000110001101011000110001101011010101100110001100111100110001100111101111011110"),
                ("1111111111110010110001100110011100111001101101101011010010000100001000010000100001000010000100001000010000100001000010000100010111101110000101000010000100001000010000100101001010010100110011100111001110011101101100111001011001110111101110010110001100"),
                ("1100111001011000110001100110011100111001100111001110011010010100101001010010100101000010000100001000010000100001000010000100010111101110000101000010000100001000010000100111000110000100110011100111011010110101101001110011110011100111001110011100111001"),
                ("1100111001011000110001100110011100111001100111001110011010010100101001010010100101000010000100001000010000100001000010000100010111101110000101000010000100001000010000100111000110000100110011100111011010110101101001110011110011100111001110011100111001"),
                ("0110001100011001100111001110011100111001110001101011010110101101001001010010100101000010000100001000010000100001000010000100010111101110000111011110110100001000010000100001001010011100011000110001001110011101101011010110110011001110011110011100111001"),
                ("1001110011110011100111001110011100111001110001101011010110101101001001010000100001000010000100001000010000100001000010000100011011110111011110111101111011101000010000100001001010010100101001010011101011010100111001110011101101011010110101101001110011"),
                ("1001110011110011100111001110011100111001110001101011010110101101001001010000100001000010000100001000010000100001000010000100011011110111011110111101111011101000010000100001001010010100101001010011101011010100111001110011101101011010110101101001110011"),
                ("1011010110100111100111001110011101011010110101001110011110101101001001010000100001000010000100001000010000100010111101111011110111101110100001000010000100001000010000100001000010000100001000010000100101001110101011010110101101001110011101100110001100"),
                ("1011010110101101011010110100111101011010100111001110011110101101001001010000100001000010000100001000101111011100001000010000100001000011101101000010000100001001010010100101001010010100001000010001100011000100111101011010110101100011000110100110001100"),
                ("1011010110101101011010110100111101011010100111001110011110101101001001010000100001000010000100001000101111011100001000010000100001000011101101000010000100001001010010100101001010010100001000010001100011000100111101011010110101100011000110100110001100"),
                ("1001110011100111101011010110101101011010101101101011010010010100101000010000100001000010000100001000101111011100001000010000110111101110000110111101110100001000010000100001000010000100101001010011101011010110100100101001010000100101001010011100011000"),
                ("1001110011100111101011010110101101011010101101101011010010010100101000010000100001000010000100001000101111011100001000010000110111101110000110111101110100001000010000100001000010000100101001010011101011010110100100101001010000100101001010011100011000"),
                ("0100101001010010100001000010001100011000100111100011000010010100101000010000100001000010000100001000101111011100001101111011101000010001101110111101110100001000010000100001000010000100111010110100100101001010010100101001010011100011000010010100001000"),
                ("0100101001010000100001000010000100101001110000100001000010000100001000010000100001000010000100001000110111101111011010000100001000010000100010111101110100001000010000100001000010001101011010110101100011000110000100101001110001100011000110000100001000"),
                ("0100101001010000100001000010000100101001110000100001000010000100001000010000100001000010000100001000110111101111011010000100001000010000100010111101110100001000010000100001000010001101011010110101100011000110000100101001110001100011000110000100001000"),
                ("0100001000010000100001000010000100001000010010100001000010000100001000010000100001000010000100001000010000100001000101111011111011110111011110111101110100001000010000100001000010001100001001010010100101001010010100101001010010100101001010010100101001"),
                ("0100001000010000100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100000001000010000110111101110100011011110110100001000010000100001000010000100101000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100000001000010000110111101110100011011110110100001000010000100001000010000100101000010000100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100011011000010000110111101111101110111101111101101000010000100001001010010100001000010000100001000010000100001000010000100101001110000100001000"),
                ("0100001000010000100001000010000100001000101111101111011010000100001000010000100001000010000100001000010000100001000010000100000001000011011110111101111101101000010000100001000010000100011011110111011110111010000100001000010001100011000100110100001000"),
                ("0100001000010000100001000010000100001000101111101111011010000100001000010000100001000010000100001000010000100001000010000100000001000011011110111101111101101000010000100001000010000100011011110111011110111010000100001000010001100011000100110100001000"),
                ("0100001000010000100001000010001101111011000011101111011010000100001000010000100001000010000100001000010000100011011101111011100001000010000111011110110100001000010000100001000010000100011011110111101111011110111101111011110110100001000010000100001000"),
                ("0100001000010000100001000010001101111011110111011110111101111011101000010000100001000010000100001000101111011110111000010000100001000010000110111101110100001000010000100001000010000100001000010001011110111101111011110111101110100001000010000100001000"),
                ("0100001000010000100001000010001101111011110111011110111101111011101000010000100001000010000100001000101111011110111000010000100001000010000110111101110100001000010000100001000010000100001000010001011110111101111011110111101110100001000010000100001000"),
                ("0100001000010000100001000010000100001000010001011110111101111011110111010000100001000010000100011011101111011101000101111011100001000010000100001000011101101000010000100001000010000100001000010001011110111101110000100001101110100001000010000100001000"),
                ("0100001000010000100001000010000100001000010001011110111101111011110111010000100001000010000100011011101111011101000101111011100001000010000100001000011101101000010000100001000010000100001000010001011110111101110000100001101110100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000110111101110111110111101110111101110000110111101110000101000010000100001000010000100001000010000100001000110111011110111110110100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000001101111011101000110111101110111101111011101000010000100001000010000100001000010000100001000010000100001000101111011110111110110100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100000001101111011101000110111101110111101111011101000010000100001000010000100001000010000100001000010000100001000101111011110111110110100001000010000100001000"),
                ("0100001000010010100101001010000100001000010000100001000010000100001000010000100001001110111101100001010000100001000101111011111011110111011101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010000100001000"),
                ("0100001000010011101011010010010100001000010000100001000010000100001001010010100101001110111101110111110111101111011110111101101000010000100011011110110100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010001100011"),
                ("0100001000010011101011010010010100001000010000100001000010000100001001010010100101001110111101110111110111101111011110111101101000010000100011011110110100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010001100011"),
                ("0100101001010011100011000010010100001000010000100001000010000100001001110101101001001010000100011011000010000110111010000100011011110111011101000010000100001000010000100001000010000100001000010000100001000010000100001000010010100101001010001111011110"),
                ("0100001000010011100011000010010100101001010011100011000010010100101000010010100101000010000100001000110111101110111101111011110111101110000111011110110100001000010000100001000010000100001000010000100001000010000100001000010010100101001110001111011110"),
                ("0100001000010011100011000010010100101001010011100011000010010100101000010010100101000010000100001000110111101110111101111011110111101110000111011110110100001000010000100001000010000100001000010000100001000010000100001000010010100101001110001111011110"),
                ("0100001000010000100101001010010100101001010011001110011110101101001000010000100001000010000100001000110111101100001000010000100001000011011110111101110100001000010000100001000010000100001001010010100101001010010100001000010000100001000110001111011110"),
                ("1001110011010010100001000010001100011000110101101011010010010100101001010000100001000010000100001000110111101100001000010000100001000010100001000010000100001000010000100001000010000100011000110001100011000110101101011010010000100101001011000110001100"),
                ("1001110011010010100001000010001100011000110101101011010010010100101001010000100001000010000100001000110111101100001000010000100001000010100001000010000100001000010000100001000010000100011000110001100011000110101101011010010000100101001011000110001100"),
                ("1011010110110100100001000010001001110011100111101011010010000100001001010010100101000010000100001000010000100010111110111101111011110110100001000010000100001000010000100001000010000100111000110000100101001110101101011010110101100011000110010110001100"),
                ("1011010110110100100001000010001001110011100111101011010010000100001001010010100101000010000100001000010000100010111110111101111011110110100001000010000100001000010000100001000010000100111000110000100101001110101101011010110101100011000110010110001100"),
                ("1011010110110100100001000010011011010110101101101011010010000100001001110101101001001010000100001000010000100001000110111101101000010000100001000010000100001000010000100111010110101001111010110101101011010110101101011010100111011010110110011100111001"),
                ("1100111001101101101011010100111011010110100111001110011010010100101000010010100111000010010100101000010000100010111000010000100001000011101101000010000100001000010000100011010110101001110011100111001110011110101101011010100111011010110110011100111001"),
                ("1100111001101101101011010100111011010110100111001110011010010100101000010010100111000010010100101000010000100010111000010000100001000011101101000010000100001000010000100011010110101001110011100111001110011110101101011010100111011010110110011100111001"),
                ("1001110011101101011010110100111011010110101101001110011100111001101000010010100101001010000100011011101111011100001000010000110111101110100001000010000100101000010000100011000110001001110011100111001110011110001001110011110011011010110110011110111101"),
                ("1011010110101101011010110101101011010110101101001110011100111001111010010010100101000110111101100001000010000100001000010000100001000010100001000010000100101001010010100001001010010100111010110101001110011110101001110011110011100111001110011111011110"),
                ("1011010110101101011010110101101011010110101101001110011100111001111010010010100101000110111101100001000010000100001000010000100001000010100001000010000100101001010010100001001010010100111010110101001110011110101001110011110011100111001110011111011110"),
                ("1111111111100111100111001101101011010110101101011010110100111001111010010010100101000101111011100001000010000100001110111101101000010000100001000010000100001001010011100011000110000100111010110101011010110100111011010110110010110001100011001111011110"),
                ("1111111111111110110001100110011100111001110011011010110110101101001001010000100001000101111011100001000010000100001101111011110111101111101101000010000100001000010000100111000110000100111010110101011010110101101100111001011000111001110111111111111111"),
                ("1111111111111110110001100110011100111001110011011010110110101101001001010000100001000101111011100001000010000100001101111011110111101111101101000010000100001000010000100111000110000100111010110101011010110101101100111001011000111001110111111111111111"),

                -- 5_explosion_3
                ("1111111111111111111011110111100110001100011001011010110010010100101000010000100001000110111101100001000010000100001000010000100001000011011110111101111101101000010000100101001010010100111010110101011010110100111100111001011000111001110111111111111111"),
                ("1111111111111111111011110111100110001100011001011010110010010100101000010000100001000110111101100001000010000100001000010000100001000011011110111101111101101000010000100101001010010100111010110101011010110100111100111001011000111001110111111111111111"),
                ("1111111111100111100111001110011100111001110011001110011010010100101000010000100001000010000100011011101111011110111000010000100001000010000100001000010000101000010000100001000010000100001001010011101011010110101001110011100110110001100100111001110011"),
                ("1011010110100111100111001110011001110011100110100101001010010100101000010000100001000010000100001000010000100001000000010000100001000010000110111101110100011011110110100011000110000100001000010000100101001110101101011010110101011010110101101100111001"),
                ("1011010110100111100111001110011001110011100110100101001010010100101000010000100001000010000100001000010000100001000000010000100001000010000110111101110100011011110110100011000110000100001000010000100101001110101101011010110101011010110101101100111001"),
                ("1011010110101101100111001110011001110011100110100101001010000100001000010000100001000010000100001000010000100010111000010000110111101111101101000010000100010111101110000101001010010100101001010011101011010110100100101001010011001110011100111001110011"),
                ("1001110011101101011010110100111101011010010010100101001010000100001000010000100001000010000100011011101111011110111000010000110111101111011101000010000100010111101110000110111101110100011000110001100011000110000100101001010010100101001010011101011010"),
                ("1001110011101101011010110100111101011010010010100101001010000100001000010000100001000010000100011011101111011110111000010000110111101111011101000010000100010111101110000110111101110100011000110001100011000110000100101001010010100101001010011101011010"),
                ("1001110011101101001110011110100100101001010010100101001010010100101000010000100001000101111011100001000010000100001000010000100001000010000110111101111011110111101111011101000010000100011000110000100101001010010100101001010000100001000010000100101001"),
                ("1011010110100111001110011110100100101001010010100001000010010100101001010000100011011000010000100001000010000100001000010000100001000010000100001000010000100001000010100001000010000100001001010011100011000010010100001000010000100101001010010100101001"),
                ("1011010110100111001110011110100100101001010010100001000010010100101001010000100011011000010000100001000010000100001000010000100001000010000100001000010000100001000010100001000010000100001001010011100011000010010100001000010000100101001010010100101001"),
                ("1101011010110100100101001010010100101001010000100001000010000100001000110111101100001000010000100001000010000100001000010000100001000010000100001000010000100001000010100011011110110100001001010011100011000010010100101001010010100101001110001100011000"),
                ("1101011010110100100101001010010100101001010000100001000010000100001000110111101100001000010000100001000010000100001000010000100001000010000100001000010000100001000010100011011110110100001001010011100011000010010100101001010010100101001110001100011000"),
                ("0100101001110100100101001010010100101001010000100001000010000100011011101111011111011101111011110111000010000100001000010000100001000010000100001000010000110111101111011110111101110100001001010011100011000110000100101001010010100101001010000001100011"),
                ("1001110011110100100001000010000100101001110110100001000010000100001000101111011111011010000100010111000010000100001000010000100001000010000100001000010000110111101110000100001000010100001001010011100011000010000100001000010000100001000010000111001110"),
                ("1001110011110100100001000010000100101001110110100001000010000100001000101111011111011010000100010111000010000100001000010000100001000010000100001000010000110111101110000100001000010100001001010011100011000010000100001000010000100001000010000111001110"),
                ("0100101001010000100001000010000100001000010000100001000010000100001000101111011111011010000100010111000010000100001000010000100001000010000100001000011011110111101111011100001000010100001000010000100101001010000100001000110111011110111110101100111001"),
                ("0100101001010011101111011101110100001000110111101111011101111011111011010000100011011000010000100001000010000100001000010000100001000010000110111101110100001000010000000100001000011101110111101111011110111010000100001000000010000100001101111100011000"),
                ("0100101001010011101111011101110100001000110111101111011101111011111011010000100011011000010000100001000010000100001000010000100001000010000110111101110100001000010000000100001000011101110111101111011110111010000100001000000010000100001101111100011000"),
                ("0100101001010001101111011010000100001000110111011110111000010000100001101111011110111000010000100001000010000100001000010000100001000010000100001000010100001000010000000100001000011101110111101110000100001101111011110111101110000100001101110000100001"),
                ("0100001000110111011110111010000100001000101110000100001101111011100001000010000100001000010000100001000010000100001000010000100001000010000110111101110100011011110111101100001000011011111011110110000100001000011101111011010001101111011101110000100001"),
                ("0100001000110111011110111010000100001000101110000100001101111011100001000010000100001000010000100001000010000100001000010000100001000010000110111101110100011011110111101100001000011011111011110110000100001000011101111011010001101111011101110000100001"),
                ("0100001000101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000101000010000000100001000011011110111110110100001000110110000100001"),
                ("0000100001000011011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111011110110000100001000010000100001101110100001000110110001100011"),
                ("0000100001000011011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000111011110110000100001000010000100001101110100001000110110001100011"),
                ("1011110111000011011110111101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111101110110001100"),
                ("1011110111000011011110111101110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111101110110001100"),
                ("0100001000110110000100001101111011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010001100011"),
                ("0100001000010001101111011101110000100001000010000100001101111011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111000010000100001000010000100001"),
                ("0100001000010001101111011101110000100001000010000100001101111011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111000010000100001000010000100001"),
                ("0100001000010001011110111101111011110111110111011110111101111011101000000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111110111101111011110111011110111000010000100001"),
                ("1101111011010000100001000010000100001000101110000100001101111011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111101111101110111101111011110111101110100001000010000100001000110111011110111"),
                ("1101111011010000100001000010000100001000101110000100001101111011110111000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000011011110111101111101110111101111011110111101110100001000010000100001000110111011110111"),
                ("0100001000010000100001000010000100001000101111011110111010000100010111101111011100001000010000100001110111101110111000010000100001000010000100001000010000100001000010100001000010000100010111101111011110111110110100001000010000100001000010000100001000"),
                ("0100001000010000100001000010000100001000010001010110101010010100111011101111011110111101111011111011000010000100001000010000100001000010000100001000010000110111101111101110111101110100010111101111011110111010000100001000010000100001000010000100001000"),
                ("0100001000010000100001000010000100001000010001010110101010010100111011101111011110111101111011111011000010000100001000010000100001000010000100001000010000110111101111101110111101110100010111101111011110111010000100001000010000100001000010000100001000"),
                ("0100101001010000100001000010010100001000010000100001000010010100101000010000100001000010000100010111000010000100001000010000100001000010000100001000011011101000010001011110111101110100001000010000100001000010000100001000010000100001000010011111011110"),
                ("1100011000110000100101001010000100101001010010100101001010000100001000010000100001000110111101110111000010000100001101111011111011110110100010111101110000100001000010000111011110110100001000010000100001000010000100001000010010100101001010000100101001"),
                ("1100011000110000100101001010000100101001010010100101001010000100001000010000100001000110111101110111000010000100001101111011111011110110100010111101110000100001000010000111011110110100001000010000100001000010000100001000010010100101001010000100101001"),
                ("0100101001010010100101001010011101011010100111100011000010010100101000010000100010111101111011110111101111011110111101111011111011110110100010111101110000100001000010000110111101110100001000010000100001000010000100101001010011100011000010000100001000"),
                ("0100101001010010100101001010011101011010100111100011000010010100101000010000100010111101111011110111101111011110111101111011111011110110100010111101110000100001000010000110111101110100001000010000100001000010000100101001010011100011000010000100001000"),
                ("0100101001010010100101001010011001110011100111100011000010010100101000010000100010111010000100010111000010000111011010000100001000010000100010111101110000110111101111011101000010000100101001010010100001000010000100101001010010100101001100111101011010"),
                ("1100011000110001100011000110101011010110100110100101001010000100001000010000100001000010000100010111000010000100001101111011110111101111011110111101110000110111101110100001000010001101011000110000100101001010010100101001110001001110011100111001110011"),
                ("1100011000110001100011000110101011010110100110100101001010000100001000010000100001000010000100010111000010000100001101111011110111101111011110111101110000110111101110100001000010001101011000110000100101001010010100101001110001001110011100111001110011"),
                ("1100111001011001001110011110100100101001110101101011010010000100001000010000100001000010000100010111000010000100001000010000100001000011011110111101110000110111101110100001000010000100101000010000100101001110101100011000100111001110011110011100111001"),
                ("1111011110111101001110011010010100101001010010100101001010010100101001010010100101000110111101100001000010000100001000010000100001000011011100001000011011110111101110100001000010000100001000010000100101001010010100101001110101100111001110011110111101"),
                ("1111011110111101001110011010010100101001010010100101001010010100101001010010100101000110111101100001000010000100001000010000100001000011011100001000011011110111101110100001000010000100001000010000100101001010010100101001110101100111001110011110111101"),
                ("1111111111111011100111001100110100101001010010100001000010010100101001010000100010111000010000100001000010000100001000010000100001000010000100001000011011110111101110100001000010000100001001010011100011000010011101011010100111100111001110011111111111"),
                ("1111111111111111100111001100110100001000010000100001000010010100101000101111011100001000010000100001000010000100001000010000100001000010000100001000010000100001000011101101000010000100001001010010100101001100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001100110100001000010000100001000010010100101000101111011100001000010000100001000010000100001000010000100001000010000100001000010000100001000011101101000010000100001001010010100101001100111100111001110011100111001111111111111111"),

                -- 6_explosion_0_0
                ("1111111111111111111111111111111111111111111111111011110011000110011001101101011010011010010100101001110001100001001010010100101001010010100011010110101001110110101101100110110101101001111001110011100111001110011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110011000110011001101101011010011010010100101001110001100001001010010100101001010010100011010110101001110110101101100110110101101001111001110011100111001110011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001101101011010011110001100001001010010100101001010010100101001010010100111000110001001110110101101100110011100111001111001110011100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110110101101011010110100111001111010100111001111010110001100001001010010100111010110101011010110101101001110110101101001111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110110101101011010110100111001111010100111001111010110001100001001010010100111010110101011010110101101001110110101101001111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110110100111001110011101101011010110101101011010110110001100011010110101100010011100111001110110101101001111001110011001110110101101100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100110110100111001111010110101101011010110101101010110010010100101001010011001110011100111001110110101101100111001110011100111001110011100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100110110100111001111010110101101011010110101101010110010010100101001010011001110011100111001110110101101100111001110011100111001110011100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001001110011101101011010110101101011010011100111001110011110001100011010010000100001001010011001110011100111011010110101101001111001110011100111001110011100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001001110011101101011010011101101011010110101101011010110110101101001000010000100001000010000100110011100111011010110101101100111001110011100111001110011100111001110011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001001110011101101011010011101101011010110101101011010110110101101001000010000100001000010000100110011100111011010110101101100111001110011100111001110011100111001110011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001011010110110011100111001101101011010110101101011010011010010100101000010000100001001010011101010110101101001110011100111100110011100111001111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001011010110110011100111001101101011010110101101011010011010010100101000010000100001001010011101010110101101001110011100111100110011100111001111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001100111001110011100110011101101011010110101101011011010010010100101001010010100111000110001001110110101101001110011100111100110110101101001111001110011111011110111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011001110011101101011010110101101011010110100111001110011100111001101001010010100101001010011001110110101101001110110101101011010011100111100111001110010110001100111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011001110011101101011010110101101011010110100111001110011100111001101001010010100101001010011001110110101101001110110101101011010011100111100111001110010110001100111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111011010110110011100111001110011100110110101101011010011010010100111000110101101011000010010100101000010001101010011100111001110110101101011010011100110110011001110011100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110011101101011011010010010100101001110101101011010110101101001001010010100111000110001001111001110011001110011100111100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110011101101011011010010010100101001110101101011010110101101001001010010100111000110001001111001110011001110011100111100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011011010110101101011010011100111001110011010010100111000010010100111000110101101001001010010100101001010011101010110101101100111001110011011010110101101011010110100111001110011111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110110101101011010011100111001110011100111001111010010010100101001010010100111000110001001110110101101001111001110011011010110101101011010110110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110110101101011010011100111001110011100111001111010010010100101001010010100111000110001001110110101101001111001110011011010110101101011010110110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110110011100111001110011100110011101101011010110100111001110011110101101011000010010100101001010010100101001010011001110110101101011011001110011001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001101101011010110101101011010110110001100001001010010100101001010010100101001010010100110110101101001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001101101011010110101101011010110110001100001001010010100101001010010100101001010010100110110101101001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001100111001110011100111001111010110001100001001110001100011000110001100001001010010100010011100111011011001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001100111001110011100111001111010110001100001001110001100011000110001100001001010010100010011100111011011001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100111001110011100101001010010100101001010010100101001010011100001000010000100110011100111100111001110011100111001110010110001100110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001110011100111001101101011010011110101101011000010010100101001010010100101001010010100111010110101001111001110011100111001110010110001100011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001110011100111001101101011010011110101101011000010010100101001010010100101001010010100111010110101001111001110011100111001110010110001100011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110011001100111001110011100110011101101011010011110101101010011101101011011000010010100101001010010100111000110000100111010110101011010011100111100111001110010110001100011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110011001100111001110011100110110101101011010011110101101010011101101011011000010010100111000110001100001001010011001110110101101001110011100111001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110011001100111001110011100110110101101011010011110101101010011101101011011000010010100111000110001100001001010011001110110101101001110011100111001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110110011100111001100111001110110101101011010011110101101010011101101011011000110101101010011100111101011010110101011010110101101011011001110011001111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110110101101011010110100111001110011100111001101001110101101010011100111101010110101101011010110101101011010011100111100111001110011100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110110101101011010110100111001110011100111001101001110101101010011100111101010110101101011010110101101011010011100111100111001110011100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100111010110001100110011100110011101101011010110100111001110110110101101001000010010100111010110101001110011100111011010110101101011011001110011100111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001001110011110011100111001100111001110110101101011010011110001100001001010010100101001010010100111000110001001110110101101011011001110011100111001110010110001100111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001001110011110011100111001100111001110110101101011010011110001100001001010010100101001010010100111000110001001110110101101011011001110011100111001110010110001100111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011001110011110011100111001110011100110110101101011010011110101101011010110001100001001010010100001001010011011010110101101011011001110011100111001110011111011110011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011001110011110011100111001110011100110110101101011010011110101101011010110001100001001010010100001001010011011010110101101011011001110011100111001110011111011110011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101110011001110011100111001111001110011100110110101101011010110101101011011010010010100101001010010100001000010001001110011100111011011001110011100111001110010110001100110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110011100111001110110101101011010011110101101001001110101101001001010010100101001010011101010110101101011010011100111100110011100111100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001100111001110011100111001110110101101011010011110101101001001110101101001001010010100101001010011101010110101101011010011100111100110011100111100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001100111001110110101101011010110101101011010011010010100111010100111001111010110100100111000110001001110110101101011011001110011100110110101101001110011110011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110110101101011010110101101011010110110101101011010100111001110011100110100111000110001001110011100111001111001110011100110110101101011010110110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110110101101011010110101101011010110110101101011010100111001110011100110100111000110001001110011100111001111001110011100110110101101011010110110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110011101101011010011100111001110110100111001110011100111001111000110001100010011100111011010110101101011011001110011100110110101101011010110110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111011001100111001110011100111001110011100110110101101011011010010010100110011100111001111010110101101010011100111001110011100111001110011100111001111001110011100111001110011001110011110011100111001110011111111111111111111111111"),
                ("1111111111111111111111111011001100111001110011100111001110011100110110101101011011010010010100110011100111001111010110101101010011100111001110011100111001110011100111001111001110011100111001110011001110011110011100111001110011111111111111111111111111"),

                -- 6_explosion_0_1
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0110001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001110010110001100111011111111111111111111101100011000110011110111101111011110011000110011111111111111101100011001111011001110011100111001110011011011111111111111101110011100111001110011100110001100011000110001100111111111111111"),
                ("1100111001110011100111001110010110001100111011111111111111111111101100011000110011110111101111011110011000110011111111111111101100011001111011001110011100111001110011011011111111111111101110011100111001110011100110001100011000110001100111111111111111"),
                ("1100111001110011100111001110011100111001110011100111001011000110011101110011100111001011000110001100110011100111001110011100111001110011100111001110011100111001110011100111001110010110001100011000110001100011001100111001110011100111001110011111111111"),
                ("1100111001110011100111001110011100111001100111001110011100111001101100110011100111001110011100111001110011100111001110011100111001110011100111001110011011011001110011100110011100111100110110101101001110011100111100111001110011100111001110011111011110"),
                ("1100111001110011100111001110011100111001100111001110011100111001101100110011100111001110011100111001110011100111001110011100111001110011100111001110011011011001110011100110011100111100110110101101001110011100111100111001110011100111001110011111011110"),
                ("1100111001110011100111001100111001110011100111100111001110011100111001100111001110011110011100111001110011100111001110011100111001110011100111001110011011011001110011100110110101101100111001110011011010110101101100111001100111001110011110010110001100"),
                ("1100111001110011100111001100111001110011100111100111001110011100111001100111001110011110011100111001110011100111001110011100111001110011100111001110011011011001110011100110110101101100111001110011011010110101101100111001100111001110011110010110001100"),
                ("1011010110100111011010110101101001110011110011100111001110011100110011101101011010110101101011010011110011100111001110011100111001110011001110110101101001110011100111011010110101101001111001110011001110011101101011010110101101011010110110011100111001"),
                ("1011010110101101011010110101101001110011110011100111001100111001110110101101011010110101101011010110110011100111001100111001110110101101011010110101101001110110101101011010110101101011010110101101011010110101101001110011100111011010110101101011010110"),
                ("1011010110101101011010110101101001110011110011100111001100111001110110101101011010110101101011010110110011100111001100111001110110101101011010110101101001110110101101011010110101101011010110101101011010110101101001110011100111011010110101101011010110"),
                ("1101011010100111011010110101101011010110101101011010110101101011010110101101011010011100111001110011110011100111001100111001110110101101011010011100111001111010110101001110110101101011010110101101011010110100111101011010100111011010110100111001110011"),
                ("0100101001100111011010110101101011010110101101011010110101101011010011100111001111010110101101011010101101011011001100111001110110101101001110011100110100101001010010100110011100111011010110101101011010110100111101011010101101001110011110000100101001"),
                ("0100101001100111011010110101101011010110101101011010110101101011010011100111001111010110101101011010101101011011001100111001110110101101001110011100110100101001010010100110011100111011010110101101011010110100111101011010101101001110011110000100101001"),
                ("1001110011101101011010110100111001110011101101001110011100111001110110100111001110011100111001110011100111001101001110101101010110101101001110011100111100001001010011100010011100111101010011100111011010110100111101011010101101101011010010010100101001"),
                ("1001110011100111101011010010011101011010101101101011010110001100011010100111001110110101101011010110110101101001001110001100011000110001101010011100110100111010110101101010011100110100101001010011101011010110001101011010101101001110011010011100011000"),
                ("1001110011100111101011010010011101011010101101101011010110001100011010100111001110110101101011010110110101101001001110001100011000110001101010011100110100111010110101101010011100110100101001010011101011010110001101011010101101001110011010011100011000"),
                ("1101011010100111101011010110100100101001110101101011010010010100101000010010100111000110001100011000110001100001001010010100101001010011100011010110101100011010110101100001001010010100101000010000100001000110101011010110101101101011010010010100101001"),
                ("1101011010100111001110011100111101011010010011100011000010010100101001110101101011010010010100101001010010100101001110001100001001010010100101001010011101011010110100100101001010010100101000010000100001000010000100101001110001100011000010010100101001"),
                ("1101011010100111001110011100111101011010010011100011000010010100101001110101101011010010010100101001010010100101001110001100001001010010100101001010011101011010110100100101001010010100101000010000100001000010000100101001110001100011000010010100101001"),
                ("1001110011110001001110011110100100101001010010100101001010010100111010100111001110011110001100001001010010100101001110001100001001010010100101001010010100101001010010100001001010011100001001010010100001000010010100101001110100100101001010010100101001"),
                ("1001110011110001001110011110100100101001010010100101001010010100111010100111001110011110001100001001010010100101001110001100001001010010100101001010010100101001010010100001001010011100001001010010100001000010010100101001110100100101001010010100101001"),
                ("1001110011110000100101001010010100101001010000100001000010010100110011110101101011010110001100001001010010100111000110001100001001010010100101001010010100101001010011101010011100111001111010110100100101001100111001110011110000100101001010010100001000"),
                ("1001110011100111100011000110000100101001010000100101001110001100010011101101011011010010010100111000010010100101000010010100101001010010100111000110000100111000110001001110110101101011010110101101001110011100111001110011100111101011010110001101011010"),
                ("1001110011100111100011000110000100101001010000100101001110001100010011101101011011010010010100111000010010100101000010010100101001010010100111000110000100111000110001001110110101101011010110101101001110011100111001110011100111101011010110001101011010"),
                ("1001110011101101001110011100111101011010100111011010110100111001110110101101011010110100111001101001010010100101001010000100001001010011001110011100111101010011100111001110011100111001110011100111011010110101101001110011100111011010110100111001110011"),
                ("1001110011101101001110011101101011010110100111011010110101101011010110101101011010110101101011011010110101101010011100111001110110101101011010110101101011011001110011011010110101101001110011100111011010110101101011010110101101011010110101101011010110"),
                ("1001110011101101001110011101101011010110100111011010110101101011010110101101011010110101101011011010110101101010011100111001110110101101011010110101101011011001110011011010110101101001110011100111011010110101101011010110101101011010110101101011010110"),
                ("1001110011101101001110011101101011010110101101011010110101101011010110101101011010110100111001110110100111001111001101101011010011100111011010011100111100110011100111011010110101101100111001110011100111001100111100111001100111001110011110011100111001"),
                ("1100111001110011100111001110011001110011110011100111001110011100111001100111001111001100111001110011110011100111001110011100111001110011100111001110011100110011100111001110011100111011010011100111100111001110011100111001110011011010110100111011010110"),
                ("1100111001110011100111001110011001110011110011100111001110011100111001100111001111001100111001110011110011100111001110011100111001110011100111001110011100110011100111001110011100111011010011100111100111001110011100111001110011011010110100111011010110"),
                ("1100111001110011100111001110011100111001110011100111001110011100111001110011100110011100111001111001110011100111001110011100111001110011001110110101101011011001110010110011001110011001110011100111100111001110011100111001100111001110011100111001110011"),
                ("1100111001101101011010110101101001110011110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110110101101011011001110011100111001110011100111001110011100111001110011100111001101101100111001110011100111001"),
                ("1100111001101101011010110101101001110011110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110110101101011011001110011100111001110011100111001110011100111001110011100111001101101100111001110011100111001"),
                ("1001110011101101011010110100111100111001011001111011110011000110011001110011100111001110011100101100011000110001100110011100111001110011100110110101101011011001110011100101100011001111011001110011100111001110011100111001110011100111001110011100111001"),
                ("1001110011101101011010110100111100111001011001111011110011000110011001110011100111001110011100101100011000110001100110011100111001110011100110110101101011011001110011100101100011001111011001110011100111001110011100111001110011100111001110011100111001"),
                ("1100111001110011100111001110010110001100110010110001100111101111001100011000110011001110011100101100011000110011001110011100111001110011100111001110011001111001110010110011110111101111001100011001100111001011000110001100011000110001100011001100111001"),
                ("1100111001110010110001100111101111011110110011111111111111111111101110111101111001100110011100111111111111111101100110011100111001110011100111001110011001111001110011111011111111111111101110011101111011110011000110001100111111111111111111101111011110"),
                ("1100111001110010110001100111101111011110110011111111111111111111101110111101111001100110011100111111111111111101100110011100111001110011100111001110011001111001110011111011111111111111101110011101111011110011000110001100111111111111111111101111011110"),
                ("1100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 6_explosion_1_0
                ("1111111111111111111011110011001100111001100111001110011100111001110110100111001111000010010100111000100111001110011110101101011010110101101001001010010100101001010011101011001110011100111001110011100111001110011100111001110010110001100111111111111111"),
                ("1111111111111111111011110011001100111001100111001110011100111001110110100111001111000010010100111000100111001110011110101101011010110101101001001010010100101001010011101011001110011100111001110011100111001110011100111001110010110001100111111111111111"),
                ("1111111111111111100111001110011001110011101101011010110101101011010110100111001101001010010100101001110101101010011010010100101001010010100101000010000100001001010010100111010110101011010011100111001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001110011001110011101101011010110110101101001001110001100001000010000100001000010000100001001010010100001000010000100001001010011100011000110001101010011100111011010110101101100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001110011001110011101101011010110110101101001001110001100001000010000100001000010000100001001010010100001000010000100001001010011100011000110001101010011100111011010110101101100111001110011100111001111111111111111"),
                ("1111111111111110110001100011001100111001110011100111001101101011010110100111001101001010010100101000010000100001000010010100101000010000100001000010000100001001010011100010011100111001111010110101001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111111111111110011100111001110011100111001101101011010110101101011010011010010100101000010000100001001010010100101001010010100101001010010100101000010001100010011100111001111010110101001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111111111111110011100111001110011100111001101101011010110101101011010011010010100101000010000100001001010010100101001010010100101001010010100101000010001100010011100111001111010110101001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111111111111111010110001100110011001110011101101011010110100111001111010010010100101000010000100001000010010100101001010010100101000010000100001000010001101010011100111101011010110101100111001110011100111001110010110001100111111111111111"),
                ("1111111111111111111011110111100110001100011001001110011100111001111010010010100101001010010100101001010000100001000010000100001000010000100001000010000100101001010011101011010110101100011010110101011010110110011100111001011000110001100111111111111111"),
                ("1111111111111111111011110111100110001100011001001110011100111001111010010010100101001010010100101001010000100001000010000100001000010000100001000010000100101001010011101011010110101100011010110101011010110110011100111001011000110001100111111111111111"),
                ("1111111111111110111001110011001001110011110011001110011110001100001001010010100111000010010100101001010010100101001010000100001000010000100111010110101100001001010011101010011100111101011010110101011010110101101100111001111010111001110111111111111111"),
                ("1111111111111110111001110011001001110011110011001110011110001100001001010010100111000010010100101001010010100101001010000100001000010000100111010110101100001001010011101010011100111101011010110101011010110101101100111001111010111001110111111111111111"),
                ("1111111111111111111111111011001011010110101101001110011010010100101001010010100111000010010100101000010000100001000010000100001000010000100111000110000100101001010011101011010110101101010011100111001110011100111100111001011001111111111111111111111111"),
                ("1111111111111111111111111011001001110011101101011010110110001100001001110001100011000010010100101000010000100001000010000100001001010011100001001010010100101001010010100101001010011101010011100111011010110101101011010110110011111111111111111111111111"),
                ("1111111111111111111111111011001001110011101101011010110110001100001001110001100011000010010100101000010000100001000010000100001001010011100001001010010100101001010010100101001010011101010011100111011010110101101011010110110011111111111111111111111111"),
                ("1111111111111110111001110011001100111001101101011010110110101101001001110101101011000010010100101001010000100001000010010100101001010010100101001010010100101001010010100101001010010100111010110101011010110101101011010110100111100111001111111111111111"),
                ("1111111111111111110111101110011100111001100111001110011110101101011010100111001111010010010100101001010000100001000010000100001001010010100101001010010100101001010010100111000110001001110110101101011010110100111001110011100111100111001111111111111111"),
                ("1111111111111111110111101110011100111001100111001110011110101101011010100111001111010010010100101001010000100001000010000100001001010010100101001010010100101001010010100111000110001001110110101101011010110100111001110011100111100111001111111111111111"),
                ("1111111111111111100111001110011011010110100111101011010100111001110110101101011011010010000100001000010000100001000010000100001001010010100101001010011100011000110000100111010110101001111010110101001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111111011110111101100111001101101011010110100111001110011100111001111010010010100101000010000100001000010000100001000010000100101001010011101011000110000100101001010010100101001010011001110011101101011010110110011110111101111111111111111"),
                ("1111111111111111111011110111101100111001101101011010110100111001110011100111001111010010010100101000010000100001000010000100001000010000100101001010011101011000110000100101001010010100101001010011001110011101101011010110110011110111101111111111111111"),
                ("1111111111111111111011110111101100111001110011011010110101101011010011100111001111010110101101011000010010100101000010000100001000010000100001000010000100101001010010100101001010010100111000110001011010110101101001110011110010110001100111111111111111"),
                ("1111111111111111110111101011001100111001100111100111001101101011010011110101101011010110001100001001010010100101000010000100001000010000100001001010010100101001010010100101001010010100111000110001001110011110011100111001110010110001100111111111111111"),
                ("1111111111111111110111101011001100111001100111100111001101101011010011110101101011010110001100001001010010100101000010000100001000010000100001001010010100101001010010100101001010010100111000110001001110011110011100111001110010110001100111111111111111"),
                ("1111111111111110111001110011001100111001100111011010110101101011010110101101011010011110001100001001010000100001000010000100001000010000100001000010000100111000110000100101001010011101011000110001001110011101101100111001110011100111001111111111111111"),
                ("1111111111111110111001110011001100111001100111011010110101101011010110101101011010011110001100001001010000100001000010000100001000010000100001000010000100111000110000100101001010011101011000110001001110011101101100111001110011100111001111111111111111"),
                ("1111111111111111110111101110011100111001110011100111001100111001110011100111001110110110101101001001010010100101000010000100001000010000100001000010000100101001010010100101001010011001110011100111001110011101101011010110110011100111001111111111111111"),
                ("1111111111111110110001100110011100111001110011100111001100111001111010100111001110011110101101001001010010100101000010010100101000010000100001001010010100101001010010100101001010011001110110101101011010110100111011010110110011100111001111111111111111"),
                ("1111111111111110110001100110011100111001110011100111001100111001111010100111001110011110101101001001010010100101000010010100101000010000100001001010010100101001010010100101001010011001110110101101011010110100111011010110110011100111001111111111111111"),
                ("1111111111111111100111001110010110001100110011001110011101101011010011110101101011010010010100111000010010100101000010000100001000010000100001000010000100001001010010100101001010011101010011100111001110011100111011010110100111100111001111111111111111"),
                ("1111111111111111111111111011000110001100100111011010110101101011010011110101101001001010010100111000010000100001000010000100001000010000100001000010000100001001010011101011010110101101011000110001101011010101101011010110100111100111001111111111111111"),
                ("1111111111111111111111111011000110001100100111011010110101101011010011110101101001001010010100111000010000100001000010000100001000010000100001000010000100001001010011101011010110101101011000110001101011010101101011010110100111100111001111111111111111"),
                ("1111111111111111111111111111011100111001101101001110011100111001110011010010100101001110001100001001010010100101000010000100001000010000100011000110000100111000110001101011010110101001111000110001101011010101101011010110100111100111001111111111111111"),
                ("1111111111111111111011110111100110001100110011001110011110001100001001010010100111000010010100101001110101101001001010000100001000010000100011000110000100101001010011101010011100111101010011100111100111001110011100111001110011100111001111111111111111"),
                ("1111111111111111111011110111100110001100110011001110011110001100001001010010100111000010010100101001110101101001001010000100001000010000100011000110000100101001010011101010011100111101010011100111100111001110011100111001110011100111001111111111111111"),
                ("1111111111111110110001100011001111011110011001011010110110101101001001010010100101001010010100101001010010100101001010000100001000010000100001001010010100101001010010100101001010011101010110101101100111001110011100111001110011100111001111111111111111"),
                ("1111111111111111111111111011100110001100110011001110011110101101010011110101101001001010000100001000010000100001000010000100001000010000100001001010011100001001010010100101001010011101010110101101011010110110011100111001110011111111111111111111111111"),
                ("1111111111111111111111111011100110001100110011001110011110101101010011110101101001001010000100001000010000100001000010000100001000010000100001001010011100001001010010100101001010011101010110101101011010110110011100111001110011111111111111111111111111"),
                ("1111111111111111111111111011100110001100110011001110011010010100110011101101011011010010010100101001010000100001000010010100101001010010100001001010011100001001010011001110011100111001110110101101001110011110011100111001011001111111111111111111111111"),
                ("1111111111111111111111111011100110001100110011001110011010010100110011101101011011010010010100101001010000100001000010010100101001010010100001001010011100001001010011001110011100111001110110101101001110011110011100111001011001111111111111111111111111"),
                ("1111111111111111001110011011100110001100100111011010110010010100111010101101011010011010010100101001010000100001000010010100101001010010100111000110000100111000110001011010011100111101010110101101011010110110010110001100011101111011110111111111111111"),
                ("1111111111111110110001100011001100111001101101001110011010010100110011101101011010011110101101001001010000100001000010000100001000010000100001001010010100111000110001101011000110001100010011100111011010110101101100111001011000110001100111111111111111"),
                ("1111111111111110110001100011001100111001101101001110011010010100110011101101011010011110101101001001010000100001000010000100001000010000100001001010010100111000110001101011000110001100010011100111011010110101101100111001011000110001100111111111111111"),
                ("1111111111111111110111101110011011010110100111001110011101101011010110100111001111000110101101001000010000100001000010000100001000010000100001000010000100001001010011100001001010011101010011100111100111001100111011010110110011100111001111111111111111"),
                ("1111111111111111100111001100111011010110101101011010110100111001110011110101101001001010010100101001010000100001000010000100001000010000100001000010000100001001010010100101001010011100010011100111100111001110011100111001110011100111001111111111111111"),
                ("1111111111111111100111001100111011010110101101011010110100111001110011110101101001001010010100101001010000100001000010000100001000010000100001000010000100001001010010100101001010011100010011100111100111001110011100111001110011100111001111111111111111"),
                ("1111111111111111100111001100111100111001110011001110011100111001111010010010100101001010000100001001010000100001000010000100001000010000100001000010000100101001010011100001001010011101010110101101011010110101101001110011110010110001100111111111111111"),
                ("1111011110011001100111001110011100111001100111100011000110001100001001010010100101000010000100001000010000100001000010000100001000010000100001001010010100111000110000100101001010011001110110101101011010110101101011010110100110110001100111111111111111"),
                ("1111011110011001100111001110011100111001100111100011000110001100001001010010100101000010000100001000010000100001000010000100001000010000100001001010010100111000110000100101001010011001110110101101011010110101101011010110100110110001100111111111111111"),

                -- 6_explosion_1_1
                ("1111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0110001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001111010110001100100111111111111111111111101100111101111011111111111111111001011000110011101011100111011101111011111011110111101100111101111010111011111111111111101110011101111011110111111111111111011001100111001110011111011110"),
                ("1100111001110011100111001111010110001100100111111111111111111111101100111101111011111111111111111001011000110011101011100111011101111011111011110111101100111101111010111011111111111111101110011101111011110111111111111111011001100111001110011111011110"),
                ("1100111001100111001110011110010110001100011100111001110011100111001100111101111011101011000110011001110011100111001011000110001100011001111011110111101100111001110010110001100011000110001100011001111011110111011100111001011001100111001110010110001100"),
                ("1100111001110011011010110101101100111001011000110001100011000110011110011000110011001011000110001100110011100111001110011100111001110011100111001110011011011001110011100110011100111011010011100110110001100011001100111001110011100111001100111100111001"),
                ("1100111001110011011010110101101100111001011000110001100011000110011110011000110011001011000110001100110011100111001110011100111001110011100111001110011011011001110011100110011100111011010011100110110001100011001100111001110011100111001100111100111001"),
                ("1001110011110011011010110100111011010110100111100111001110011100101100110011100110110100111001111001110011100111001100111001110011100111100110110101101001110011100111011010110101101011011001110010110001100110011100111001110011100111001101101001110011"),
                ("1100011000100111011010110100111001110011101101001110011100111001110110100111001110011101101011010011110011100111001101101011011001110011011010110101101101010011100111011010110101101001110011100111001110011100111100111001110011001110011101101001110011"),
                ("1100011000100111011010110100111001110011101101001110011100111001110110100111001110011101101011010011110011100111001101101011011001110011011010110101101101010011100111011010110101101001110011100111001110011100111100111001110011001110011101101001110011"),
                ("1100011000100111001110011101100100101001010010100101001110101101011010110001100010011101101011010110100111001110011101101011010110101101011010011100111001111010110101101011000110000100111000110001001110011101101011010110101101011010110101101001110011"),
                ("1100011000100111001110011101100100101001010010100101001110101101011010110001100010011101101011010110100111001110011101101011010110101101011010011100111001111010110101101011000110000100111000110001001110011101101011010110101101011010110101101001110011"),
                ("0100101001110101001110011101101001110011110101001110011100111001101001010010100110011100111001110011110101101010011101101011010011100111001110011100111011011010110100100101001010010100101001010011101011010101101011010110101101011010110101101011010110"),
                ("0100101001010011101011010100111011010110101101011010110110101101001001010010100101001110101101011010100111001110011101101011011010110101001110011100111011010011100111101011000110000100101001010010100101001100111011010110100111101011010100111001110011"),
                ("0100101001010011101011010100111011010110101101011010110110101101001001010010100101001110101101011010100111001110011101101011011010110101001110011100111011010011100111101011000110000100101001010010100101001100111011010110100111101011010100111001110011"),
                ("0100001000010010100101001110001001110011100111101011010010010100101001110001100001001010010100111010100111001110110100111001111010110101101011010110101101011010110101100011000110001100011000110000100101001110101001110011010010100101001010011100011000"),
                ("0100001000010000100101001110101101011010010010100101001010000100001001010010100111000010010100101001110101101011010110001100011000110001101001001010010100001001010010100101001010010100101001010010100101001010010100101001010011100011000010010100101001"),
                ("0100001000010000100101001110101101011010010010100101001010000100001001010010100111000010010100101001110101101011010110001100011000110001101001001010010100001001010010100101001010010100101001010010100101001010010100101001010011100011000010010100101001"),
                ("0100001000010010100101001010000100101001010010100101001010000100001001010010100101001110001100011000010010100101001010010100101001010011100001000010000100001001010010100101000010000100001001010010100101001010000100001000010000100001000010011100011000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001001110101101001001010000100001001010010100101001010000100001001010010100101000010000100001000010000100001000010000100001001010010100001000010000100001000010000100001000110101001110011"),
                ("0100001000010000100001000010000100001000010000100001000010000100001001110101101001001010000100001001010010100101001010000100001001010010100101000010000100001000010000100001000010000100001001010010100001000010000100001000010000100001000110101001110011"),
                ("0100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100001000010000100101001010000100001000100111001110011"),
                ("0100001000010000100001000010000100001000010010100101001010000100001000010000100001000010000100001000010010100101000010000100001000010000100001000010000100001000010000100101000010000100001000010000100001000010010100101001010010100001000010011101011010"),
                ("0100001000010000100001000010000100001000010010100101001010000100001000010000100001000010000100001000010010100101000010000100001000010000100001000010000100001000010000100101000010000100001000010000100001000010010100101001010010100001000010011101011010"),
                ("0100001000010000100001000010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010010100001000010000100001000010010100101001010000100101001010011101011010"),
                ("0100001000010000100001000010000100001000010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010010100001000010000100001000010010100101001010000100101001010011101011010"),
                ("0100001000010000100001000010000100001000010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001010010100111000110000100101001010010100001000010010100101001010000100001000010011101011010"),
                ("0100101001010000100001000010000100101001110000100101001010010100101001110001100011000010000100001000010010100101000010000100001001010010100001001010010100101001010010100101001010011100011010110100100001000010000100101001010000100001000010000100101001"),
                ("0100101001010000100001000010000100101001110000100101001010010100101001110001100011000010000100001000010010100101000010000100001001010010100001001010010100101001010010100101001010011100011010110100100001000010000100101001010000100001000010000100101001"),
                ("0100101001010010100001000010000100101001010011100011000110001100001001010010100101001010000100001000010010100101001010010100101001010010100111010110101100001001010010100101001010010100111000110000100101001010000100101001010000100001000010000100101001"),
                ("1100011000010010100101001010011100011000110000100101001010010100101001010010100111000010010100101001010010100101001110001100001001010010100111000110001100001001010010100101001010010100101001010010100101001010000100001000010010100101001010010100101001"),
                ("1100011000010010100101001010011100011000110000100101001010010100101001010010100111000010010100101001010010100101001110001100001001010010100111000110001100001001010010100101001010010100101001010010100101001010000100001000010010100101001010010100101001"),
                ("0100101001110000100101001110001101011010101101001110011010010100101001110101101011010110101101001001010010100101001010010100101001010010100101001010010100101001010010100101001010011101011010110101101011010110101100011000110001100011000010011101011010"),
                ("0100101001010010100101001010011100011000100111001110011010010100101001100111001111010110101101001001010010100101001010010100101001010010100101001010011101011000110000100101001010011101010011100111101011010100111001110011100111100011000110101100111001"),
                ("0100101001010010100101001010011100011000100111001110011010010100101001100111001111010110101101001001010010100101001010010100101001010010100101001010011101011000110000100101001010011101010011100111101011010100111001110011100111100011000110101100111001"),
                ("1001110011110101100011000110101100011000110101001110011110101101011010110101101010011110101101011010100111001110011110101101001001010010100101001010011001110011100110100111010110101101011010110101100011000110101001110011100111101011010101101100111001"),
                ("1011010110101101001110011100111001110011101101011010110101101011010110100111001111000110001100010011101101011010011110001100011000110001100001001010011101010110101101101010011100111001111010110101101011010110101101011010110101001110011100111100111001"),
                ("1011010110101101001110011100111001110011101101011010110101101011010110100111001111000110001100010011101101011010011110001100011000110001100001001010011101010110101101101010011100111001111010110101101011010110101101011010110101001110011100111100111001"),
                ("1011010110101101100111001110011011010110101101001110011101101011011001110011100111010110101101010011101101011010011100111001110011100111011010011100111001110110101101011010110101101001110110101101011010110110011001110011100111011010110100111100111001"),
                ("1011010110101101100111001110011011010110101101001110011101101011011001110011100111010110101101010011101101011010011100111001110011100111011010011100111001110110101101011010110101101001110110101101011010110110011001110011100111011010110100111100111001"),
                ("1011010110101101100111001100111011010110110011100111001110011100111001110011100110110101101011010011100111001110110101101011011001110011011010110101101001110011100111011010110101101001110110101101100111001110011001110011100111011010110100111100111001"),
                ("1011010110100111100111001101101100111001011001100111001110011100111001110011100110110101101011010110101101011010110110011100111001110011001110110101101100110011100111011010110101101100111001110011100111001110011100111001110011100111001110011100111001"),
                ("1011010110100111100111001101101100111001011001100111001110011100111001110011100110110101101011010110101101011010110110011100111001110011001110110101101100110011100111011010110101101100111001110011100111001110011100111001110011100111001110011100111001"),
                ("1001110011110011100111001110010110001100011100110001100110011100111001110011100110011100111001110011110011100111001110011100111001110011100111001110011100110011100111001111001110010110011101111010110001100110011100111001110011100111001110011100111001"),
                ("0110001100011001100111001110010110001100111101111111111111111111111001110011100111001110011100111001110011100111001110011100101100011000110011101111011100111001110011100111111111111111101110011100110001100011001100111001110011100111001110010110001100"),
                ("0110001100011001100111001110010110001100111101111111111111111111111001110011100111001110011100111001110011100111001110011100101100011000110011101111011100111001110011100111111111111111101110011100110001100011001100111001110011100111001110010110001100"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 6_explosion_2_0
                ("1111111111011000110001100110011001110011101101001110011110001100001001010000100001001010000100001000110111101111011101111011111011110110100001000010000100101001010011101001001010010100111010110101001110011101101011010110101101100111001111101111111111"),
                ("1111111111011000110001100110011001110011101101001110011110001100001001010000100001001010000100001000110111101111011101111011111011110110100001000010000100101001010011101001001010010100111010110101001110011101101011010110101101100111001111101111111111"),
                ("1111111111011001100111001110011001110011101101001110011110101101010011110001100001001010000100001000010000100011011000010000110111101110100001000010000100101001010011101001001010010100111010110101101011010100111011010110101101001110011011001111111111"),
                ("1111111111110011100111001110011001110011101101011010110100111001110011110101101001001010000100001000010000100001000101111011110111101110000110111101110100001000010000100001000010000100111010110101001110011100111101011010101101100111001110011111111111"),
                ("1111111111110011100111001110011001110011101101011010110100111001110011110101101001001010000100001000010000100001000101111011110111101110000110111101110100001000010000100001000010000100111010110101001110011100111101011010101101100111001110011111111111"),
                ("1111111111011000110001100110011011010110101101011010110110101101001001110001100001000010000100001000010000100011011101111011110111101111011100001000011011101000010000100001000010000100001000010000100101001110001101011010101101100111001011001111111111"),
                ("1111111111111101110111101011001011010110101101001110011110001100001001010010100101000010000100001000010000100001000110111101110111101110000111011110110100001000010000100001000010000100001000010000100101001010011001110011101100110001100011101111111111"),
                ("1111111111111101110111101011001011010110101101001110011110001100001001010010100101000010000100001000010000100001000110111101110111101110000111011110110100001000010000100001000010000100001000010000100101001010011001110011101100110001100011101111111111"),
                ("1111111111111111111111111111101001110011101101011010110110101101001001010010100101000010000100001000010000100001000101111011110111101110000101000010000100001000010000100001000010000100111010110101001110011101101011010110101100110001100011101111111111"),
                ("1111111111111111111111111111101100111001100111011010110101101011011010010000100001000010000100001000010000100001000010000100011011110110000101000010000100001000010000100001000010000100001001010011101011010101101011010110110010110001100111111111111111"),
                ("1111111111111111111111111111101100111001100111011010110101101011011010010000100001000010000100001000010000100001000010000100011011110110000101000010000100001000010000100001000010000100001001010011101011010101101011010110110010110001100111111111111111"),
                ("1111111111011001111011110111011100111001101101011010110101101011010011010000100001000010010100101001010000100001000010000100001000010001011111011110111101101000010000100001000010001101011010110101101011010101101011010110110011111011110111111111111111"),
                ("1111111111011001111011110111011100111001101101011010110101101011010011010000100001000010010100101001010000100001000010000100001000010001011111011110111101101000010000100001000010001101011010110101101011010101101011010110110011111011110111111111111111"),
                ("1111111111010010110001100110011100111001101101011010110100111001110011110001100001000010010100101000010000100010111110111101101000010000100011011110111011101000010000100011000110001001110110101101001110011101101011010110011001111011110110011111111111"),
                ("1111111111010001001110011110011011010110101101001110011110001100001001010000100001000010010100101000010000100000001000010000100001000010000100001000011011111011110110100001000010000100111010110101001110011110101001110011011001100111001100111111111111"),
                ("1111111111010001001110011110011011010110101101001110011110001100001001010000100001000010010100101000010000100000001000010000100001000010000100001000011011111011110110100001000010000100111010110101001110011110101001110011011001100111001100111111111111"),
                ("1111111111010001100111001110011001110011100111001110011010010100101001010000100001000010000100001000010000100000001000010000100001000010000100001000010000110111101110100001000010000100001001010011101011010100111001110011110011100111001110011111111111"),
                ("1111111111010000001100011011000110001100110101001110011100111001111010010010100111000010000100001000010000100010111101111011110111101110000110111101111011111011110110100001001010010100001000010001001110011101101001110011011001100111001011001111111111"),
                ("1111111111010000001100011011000110001100110101001110011100111001111010010010100111000010000100001000010000100010111101111011110111101110000110111101111011111011110110100001001010010100001000010001001110011101101001110011011001100111001011001111111111"),
                ("1111111111010001101011010110101100111001100111101011010101101011010011110101101011000010010100101000110111101100001101111011100001000010000111011110110100001000010000100001001010010100110011100111011010110100111100111001110011100111001111101111111111"),
                ("1111111111110001100111001101101100111001100111011010110101101011010011010010100101001010010100101000010000100010111000010000110111101111011101000010000100001000010000100101000010000100110110101101011010110101101011010110110011100111001111101111111111"),
                ("1111111111110001100111001101101100111001100111011010110101101011010011010010100101001010010100101000010000100010111000010000110111101111011101000010000100001000010000100101000010000100110110101101011010110101101011010110110011100111001111101111111111"),
                ("1111111111110001100111001110011100111001110011001110011101101011010011110001100001000010000100001000010000100010111101111011111011110111101101000010000100001001010010100101000010001001110110101101001110011101101011010110110010110001100011101111111111"),
                ("1111111111010001100111001110011100111001110011100111001101101011010110110101101001000010010100101001010000100001000101111011111011110110100001000010000100001001010011100011010110101001110110101101001110011101101011010110110011100111001011001111111111"),
                ("1111111111010001100111001110011100111001110011100111001101101011010110110101101001000010010100101001010000100001000101111011111011110110100001000010000100001001010011100011010110101001110110101101001110011101101011010110110011100111001011001111111111"),
                ("1111111111110001100111001110011100111001110011100111001100111001111010010000100001000010010100101000010000100001000010000100010111101111011101000010000100001001010010100101001010011001110011100111101011010100111001110011110011100111001110011111111111"),
                ("1111111111110001100111001110011100111001110011100111001100111001111010010000100001000010010100101000010000100001000010000100010111101111011101000010000100001001010010100101001010011001110011100111101011010100111001110011110011100111001110011111111111"),
                ("1111111111110101100111001101101011010110100111001110011110101101001000010000100001001010010100101001010000100011011000010000110111101111011110111101111101101000010000100101000010000100011010110100100101001110101001110011110011100111001110011111111111"),
                ("1111111111110000110001100110011011010110100111011010110101101011001001010010100101000010000100001000010000100001000010000100010111101110000100001000011011111011110110100001001010010100001001010011001110011100111001110011110011100111001110011111111111"),
                ("1111111111110000110001100110011011010110100111011010110101101011001001010010100101000010000100001000010000100001000010000100010111101110000100001000011011111011110110100001001010010100001001010011001110011100111001110011110011100111001110011111111111"),
                ("1111111111010011110111101110011100111001100111011010110100111001111010010000100001000010000100001000010000100011011101111011110111101111101110111101111101101000010000100001000010000100011010110101011010110101101100111001110011100111001110011111111111"),
                ("1111111111011101110111101110011100111001100111011010110110101101001001010000100001000010000100001000010000100011011000010000110111101110100001000010000100001000010000100001000010000100110011100111011010110100111001110011110011100111001110011111111111"),
                ("1111111111011101110111101110011100111001100111011010110110101101001001010000100001000010000100001000010000100011011000010000110111101110100001000010000100001000010000100001000010000100110011100111011010110100111001110011110011100111001110011111111111"),
                ("1111111111111111111111111011001100111001101101011010110100111001101001010000100001000010000100001000010000100011011110111101101000010000100001000010000100001000010000100001000010000100011010110101001110011110011100111001011001011010110110011111111111"),
                ("1111111111111111111111111111101111011110110011011010110101101011011010010000100001000010000100001000010000100001000010000100001000010000100011011110111101101000010000100001001010010100110011100111101011010110001100111001111011001110011111111111111111"),
                ("1111111111111111111111111111101111011110110011011010110101101011011010010000100001000010000100001000010000100001000010000100001000010000100011011110111101101000010000100001001010010100110011100111101011010110001100111001111011001110011111111111111111"),
                ("1111111111111100110001100011000110001100100111011010110100111001110011010010100101001010010100101001010000100001000010000100010111101110000110111101110100001000010000100011000110001001110011100111101011010010011001110011011000111001110111111111111111"),
                ("1111111111111100110001100111101100111001100111011010110110101101001001010010100101001010010100101000010000100001000110111101110111101111011111011110110100001000010000100011010110101001111010110101011010110100111101011010100110110001100111011111111111"),
                ("1111111111111100110001100111101100111001100111011010110110101101001001010010100101001010010100101000010000100001000110111101110111101111011111011110110100001000010000100011010110101001111010110101011010110100111101011010100110110001100111011111111111"),
                ("1111111111110011100111001110011001110011101101001110011010010100111000010000100001000010000100001000010000100001000010000100010111101111011110111101110100001000010000100011000110001011010011100111001110011100111101011010100111100111001011001111111111"),
                ("1111111111110011100111001110011001110011101101001110011010010100111000010000100001000010000100001000010000100001000010000100010111101111011110111101110100001000010000100011000110001011010011100111001110011100111101011010100111100111001011001111111111"),
                ("1111111111100111100111001100111011010110101101001110011100111001110011010010100101000010010100101000010000100001000010000100010111101110000111011110110100001000010000100001001010011001110011100111001110011100111001110011101101011010110011001111111111"),
                ("1111111111100111011010110101101011010110101101001110011101101011010011010010100101001010000100001001010000100001000010000100010111101110000101000010000100001001010010100101001010010100101001010011001110011101101011010110101101011010110110011111111111"),
                ("1111111111100111011010110101101011010110101101001110011101101011010011010010100101001010000100001001010000100001000010000100010111101110000101000010000100001001010010100101001010010100101001010011001110011101101011010110101101011010110110011111111111"),
                ("1111111111110011001110011100111011010110100111101011010101101011011010010010100101001010000100001000010000100001000110111101100001000011011111011110110100111000110000100101001010010100101001010011001110011110011001110011110011001110011110011111111111"),
                ("1111111111111101100111001110011100111001100110100101001100111001110011100111001111010010010100101000010000100001000000010000110111101111011111011110110100001001010010100101001010010100101000010001101011010110011100111001110011100111001110011111111111"),
                ("1111111111111101100111001110011100111001100110100101001100111001110011100111001111010010010100101000010000100001000000010000110111101111011111011110110100001001010010100101001010010100101000010001101011010110011100111001110011100111001110011111111111"),
                ("1111111111111101100111001110011100111001100111001110011110101101010011101101011010011110101101001001010000100010111000010000110111101111101101000010000100001001010011100001000010000100001000010000100101001101101001110011110011100111001110011111111111"),
                ("1111111111100111011010110101101001110011101101011010110100111001110011101101011010011110001100001000010000100010111010000100001000010000100001000010000100001001010011100011000110000100101000010000100101001010010100101001110011100111001110011110111101"),
                ("1111111111100111011010110101101001110011101101011010110100111001110011101101011010011110001100001000010000100010111010000100001000010000100001000010000100001001010011100011000110000100101000010000100101001010010100101001110011100111001110011110111101"),

                -- 6_explosion_2_1
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1001110011111101111011110110011001110011100111100111001111101111011110111111111111111011100111001001110001100011010110001100001000010001100011000110000100001000010000100001000010000100101100011001111111111111111111011110011001100111001011000110001100"),
                ("1011010110110011100111001100111011010110110011100111001011000110001100111111111111111111011110111101011000110011001110011100111001110011100111001110011101000011000111100110011100110110011110111101111111111111111110111101011001100111001110010110001100"),
                ("1011010110110011100111001100111011010110110011100111001011000110001100111111111111111111011110111101011000110011001110011100111001110011100111001110011101000011000111100110011100110110011110111101111111111111111110111101011001100111001110010110001100"),
                ("1011010110110011100111001100111011010110100111100111001111101111001100111101111001100110011100111001110011100110110110011100111001110011100110110101101101001100011001100111001110011100111101111011111011110111100110001100110011100111001110011100111001"),
                ("1001110011110011100111001101101011010110101101001110011110011100101100111101111011001110011100111001101101011010110110011100111001110011100111001110011100101100011001001110110101101100111001110011100111001100111011010110101101001110011100111001110011"),
                ("1001110011110011100111001101101011010110101101001110011110011100101100111101111011001110011100111001101101011010110110011100111001110011100111001110011100101100011001001110110101101100111001110011100111001100111011010110101101001110011100111001110011"),
                ("1011010110100111001110011100111011010110101101011010110100111001110011110011100110110100111001110011100111001110011110011100111001110011100110011100111001111010110101001110110101101011010110101101001110011101101011010110101101011010110101101011010110"),
                ("1011010110100110100101001110101001110011100111001110011101101011010110101101011010110101101011010110101101011010011110011100111001110011001110110101101101010011100111001110011100111011010110101101011010110101101001110011101101011010110100111001110011"),
                ("1011010110100110100101001110101001110011100111001110011101101011010110101101011010110101101011010110101101011010011110011100111001110011001110110101101101010011100111001110011100111011010110101101011010110101101001110011101101011010110100111001110011"),
                ("1001110011110101001110011101101011010110100110100101001110101101010011101101011010011110101101010011101101011011010100111001110110101101011010110101101011010011100110100111000110001001110110101101011010110110101100011000110101001110011110101100011000"),
                ("1001110011110101001110011101101011010110100110100101001110101101010011101101011010011110101101010011101101011011010100111001110110101101011010110101101011010011100110100111000110001001110110101101011010110110101100011000110101001110011110101100011000"),
                ("1001110011100111001110011110101001110011100111100011000010010100110011110101101001001010010100111010010010100101000110101101010110101101001110011100111001111010110100100101001010011001110011100111101011010010010100101001010011001110011100110100101001"),
                ("1011010110101101001110011010010100101001010010100001000010010100101001010000100001000010000100001000010010100101000010000100011010110101100001001010011101001001010010100001000010001100001000010000100001000010010100101001110001101011010110000100001000"),
                ("1011010110101101001110011010010100101001010010100001000010010100101001010000100001000010000100001000010010100101000010000100011010110101100001001010011101001001010010100001000010001100001000010000100001000010010100101001110001101011010110000100001000"),
                ("1001110011100111101011010010010100101001010000100001000010010100101001010000100001000010000100001000010000100001001010000100001000010000100001001010011100011000110000100001000010000100001000010000100001000010000100001000010000100101001010010100101001"),
                ("1100011000110100100101001010000100001000010010100001000010010100101001010000100001000010000100001000010000100001001010010100101001010010100001001010010100101000010000100001001010010100101001010010100001000010000100001000010000100001000010000100001000"),
                ("1100011000110100100101001010000100001000010010100001000010010100101001010000100001000010000100001000010000100001001010010100101001010010100001001010010100101000010000100001001010010100101001010010100001000010000100001000010000100001000010000100001000"),
                ("0100001000010010100001000010000100101001010000100001000010000100001001010000100001000010000100001000010000100001001010000100001001010010100001000010000100001000010000100001000010000100001001010010100001000010000100001000010000100001000010000100001000"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010001101101000010000100001000010000100001000010000100001000010000100001000010000100001000010001101111011"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010001101101000010000100001000010000100001000010000100001000010000100001000010000100001000010001101111011"),
                ("1011110111101110100001000010000100001000010000100001000010000100001000010000100011011110111101111011010000100011011010000100001000010001011110111101110000110111101110000100001000011011101000010000100001000010000100001000110110100001000110111101111011"),
                ("0100001000000010000100001110110100001000010000100001000110111101101000010000100011011000010000110111010000100000001010000100010111101111011100001000011011110111101110000100001000011101101000010000100001000101111101111011101111011110111000011011110111"),
                ("0100001000000010000100001110110100001000010000100001000110111101101000010000100011011000010000110111010000100000001010000100010111101111011100001000011011110111101110000100001000011101101000010000100001000101111101111011101111011110111000011011110111"),
                ("0100001000101111011110111000011011110111101111011110111101111011110111010000100001000101111011110111101111011110111101111011111011110111101110111101110000110111101110000100001000010100001000010001101111011101111011110111101111011110111101111101111011"),
                ("0100001000101111011110111000011011110111101111011110111101111011110111010000100001000101111011110111101111011110111101111011111011110111101110111101110000110111101110000100001000010100001000010001101111011101111011110111101111011110111101111101111011"),
                ("0100001000110111011110111101110000100001000011011110111101111011100001010000100001000010000100011011000010000110111101111011101000010001101110111101110000100001000010000100001000010100010111101110000100001000010000100001101110000100001010000100001000"),
                ("0100001000010001101111011110110100001000110111011110111110111101110111110111101101000010000100010111000010000110111010000100001000010000100001000010001101110111101110000100001000011101111011110110100001000010001101111011000011011110111010000100001000"),
                ("0100001000010001101111011110110100001000110111011110111110111101110111110111101101000010000100010111000010000110111010000100001000010000100001000010001101110111101110000100001000011101111011110110100001000010001101111011000011011110111010000100001000"),
                ("0100001000010000100001000010010100001000010000100001000010000100001000110111101101000010000100011011101111011111011010000100001000010000100001000010000100010111101110000110111101111011111011110110100001000010000100001000101110100001000010010100101001"),
                ("0100101001010010100101001110000100101001010000100001000010000100001000010000100001000010000100001000110111101101000010010100101001010010100101000010000100011011110111011111011110110100001000010000100001000010000100001000010000100001000010010100101001"),
                ("0100101001010010100101001110000100101001010000100001000010000100001000010000100001000010000100001000110111101101000010010100101001010010100101000010000100011011110111011111011110110100001000010000100001000010000100001000010000100001000010010100101001"),
                ("1100011000110000100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001001010010100111000110000100101001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000110101101011010"),
                ("1100011000010000100101001010010100101001010011100011000110101101011000010010100101000010000100001000010010100101000010010100111010110100100001000010000100101001010010100001000010001100001000010000100001000010000100001000010000100001000010010100101001"),
                ("1100011000010000100101001010010100101001010011100011000110101101011000010010100101000010000100001000010010100101000010010100111010110100100001000010000100101001010010100001000010001100001000010000100001000010000100001000010000100001000010010100101001"),
                ("0100101001010000100101001010010100101001100111011010110100111001110011010010100101000010010100101000010000100001000100111001110011100111001101001010010100101000010000100001001010011001111010110100100001000010010100001000010000100101001010010100101001"),
                ("0100001000010000100001000010010100101001100111001110011110101101010011100111001111010100111001111010010010100111010100111001110110101101011010110101101001101000010000100111010110101011011010110100100101001110100100001000010001101011010110101101011010"),
                ("0100001000010000100001000010010100101001100111001110011110101101010011100111001111010100111001111010010010100111010100111001110110101101011010110101101001101000010000100111010110101011011010110100100101001110100100001000010001101011010110101101011010"),
                ("0100101001010011101011010100111001110011100111001110011101101011011010110101101010011101101011010110100111001101001110101101010011100111001110110101101011010011100111101010011100111001111010110101101011010100110100101001010011001110011110101001110011"),
                ("0100101001010011101011010100111001110011100111001110011101101011011010110101101010011101101011010110100111001101001110101101010011100111001110110101101011010011100111101010011100111001111010110101101011010100110100101001010011001110011110101001110011"),
                ("0100101001101101100111001110011011010110100111001110011100111001101001110001100011001100111001110110100111001111010100111001110110101101011010110101101001110110101101001111010110101011010110101101011010110101100100101001110001001110011100111011010110"),
                ("0100101001100111100111001100111011010110100111101011010110101101010011110011100111001100111001111001100111001110011100111001110110101101011010110101101100110011100111001110011100111011010110101101011010110101101001110011110101101011010101101011010110"),
                ("0100101001100111100111001100111011010110100111101011010110101101010011110011100111001100111001111001100111001110011100111001110110101101011010110101101100110011100111001110011100111011010110101101011010110101101001110011110101101011010101101011010110"),
                ("1100111001110011100111001110011011010110101101001110011100111001101100111011110101100110011100111001110011100111001110011100111001110011100111001110011100101100011001100101100011000110011001110011100111001101101011010110101101011010110101101011010110"),
                ("1100111001110011100111001100111011010110101101100111001011000110001110100111001110110110011100111001110011100111001110011100111001110010110011001110011100111001110011100111001110011111011110111100110001100011000110001100110011100111001100111100111001"),
                ("1100111001110011100111001100111011010110101101100111001011000110001110100111001110110110011100111001110011100111001110011100111001110010110011001110011100111001110011100111001110011111011110111100110001100011000110001100110011100111001100111100111001"),
                ("1100111001110011100111001110011100111001011000110001100111011110111111111111111111001110011100111001110011100111001110011100101100011000111011110111101111001100011001100110011100111100111111111111111111111011100111001110011001100111001011001111011110"),
                ("1111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 6_explosion_3_0
                ("1011010110100111001110011101101011010110101101011010110101101011010110100111001101001010000100001000010000100001000010000100001000010000100001000010000100001001010010100111010110100100001000010000100001000010011001110011100111100111001011000110001100"),
                ("1011010110100111001110011101101011010110101101011010110101101011010110100111001101001010000100001000010000100001000010000100001000010000100001000010000100001001010010100111010110100100001000010000100001000010011001110011100111100111001011000110001100"),
                ("0110001100110011100111001100111001110011101101001110011100111001110011110101101001001010000100011011101111011100001110111101101000010000100011011110111101101000010000100001000010000100001000010000100001000010000100101001010011001110011110011100111001"),
                ("1110111101111100110001100100111011010110100110100101001010000100001000010000100001000110111101100001000010000100001110111101101000010001011100001000011011101000010000100001000010000100101000010000100101001010010100101001110101100111001110011111111111"),
                ("1110111101111100110001100100111011010110100110100101001010000100001000010000100001000110111101100001000010000100001110111101101000010001011100001000011011101000010000100001000010000100101000010000100101001010010100101001110101100111001110011111111111"),
                ("1111111111111110110001100110011100111001100110100101001010000100001000010000100001000101011010110111000010000110111101111011110111101110000100001000011011111011110110100101001010010100101000010001100011000110101101011010100111100111001111111111111111"),
                ("1111111111111111110111101110011100111001110100100101001010010100101000010000100001000010000100001000101111011111011000010000100001000010000100001000010000110111101110100001000010000100101000010001100011000100111011010110100111100111001111111111111111"),
                ("1111111111111111110111101110011100111001110100100101001010010100101000010000100001000010000100001000101111011111011000010000100001000010000100001000010000110111101110100001000010000100101000010001100011000100111011010110100111100111001111111111111111"),
                ("1111111111111111100111001101101100111001110100100001000010010100101001010010100101001010000100001000101111011100001000010000100001000011011100001000010000100001000011101101000010000100101001010011100011000101101100111001110011100111001011001111111111"),
                ("1111111111111110110001100101101011010110100110100001000010010100101000010010100101001010010100111011101111011100001110111101110111101111011100001000010000100001000011011101000010000100001001010011100011000100111011010110100111100111001111100111001110"),
                ("1111111111111110110001100101101011010110100110100001000010010100101000010010100101001010010100111011101111011100001110111101110111101111011100001000010000100001000011011101000010000100001001010011100011000100111011010110100111100111001111100111001110"),
                ("1111111111111111001110011101101011010110100110100101001110001100001001010010100101000010000100001000000010000110111110111101100001000010000100001000011011110111101110100001000010000100001001010010100101001100111011010110101101100111001011000110001100"),
                ("1111111111111111001110011101101011010110100110100101001110001100001001010010100101000010000100001000000010000110111110111101100001000010000100001000011011110111101110100001000010000100001001010010100101001100111011010110101101100111001011000110001100"),
                ("1111111111111111011010110101101011010110100110100101001010010100111000010010100101000010000100001000110111101100001000010000110111101110000100001000011011101000010000100001000010000100001000010001101011010101101011010110101101011010110100111100111001"),
                ("0110001100101101001110011110101001110011110101100011000010010100101001010010100101000010000100011011101111011100001000010000110111101111101100001000011011101000010001101101000010000100001000010000100101001100111001110011100111100111001110011100111001"),
                ("0110001100101101001110011110101001110011110101100011000010010100101001010010100101000010000100011011101111011100001000010000110111101111101100001000011011101000010001101101000010000100001000010000100101001100111001110011100111100111001110011100111001"),
                ("1100111001100111001110011110100100101001010010100101001010000100001000010000100001000010000100010111000010000100001000010000111011110110100010111101110000100001000011011101000010000100001000010000100001000010011101011010110011100111001110011111111111"),
                ("1100111001110011011010110100110100101001010010100001000010000100001000010000100001000010000100010111000010000100001000010000100001000010000100001000011011101000010000100001000010000100001000010000100101001110101011010110101101011010110111111111111111"),
                ("1100111001110011011010110100110100101001010010100001000010000100001000010000100001000010000100010111000010000100001000010000100001000010000100001000011011101000010000100001000010000100001000010000100101001110101011010110101101011010110111111111111111"),
                ("1101011010110011011010110110100100101001110000100001000010000100001001010000100001000110111101100001000010000100001000010000110111101110000110111101110000111011110110100001000010000100001001010010100101001110101011010110101101011010110111111111111111"),
                ("1100111001110011011010110100111101011010100111100011000010010100101001010000100001000110111101100001000010000100001000010000110111101110000101000010001101111011110110100001000010000100001001010011100011000100111011010110101101011010110111111111111111"),
                ("1100111001110011011010110100111101011010100111100011000010010100101001010000100001000110111101100001000010000100001000010000110111101110000101000010001101111011110110100001000010000100001001010011100011000100111011010110101101011010110111111111111111"),
                ("1011010110110011100111001101101011010110101101101011010010000100001001010000100001000010000100011011000010000110111101111011110111101111011110111101110100001000010000100001000010000100101001010010100101001110101101011010100111011010110111111111111111"),
                ("0110001100100111100111001101101011010110100111100011000010010100101001010010100111011101111011111011101111011101000010000100001000010001101110111101111101101000010000100001000010000100101001010010100101001110101101011010100111001110011110011110111101"),
                ("0110001100100111100111001101101011010110100111100011000010010100101001010010100111011101111011111011101111011101000010000100001000010001101110111101111101101000010000100001000010000100101001010010100101001110101101011010100111001110011110011110111101"),
                ("1100111001100111011010110100111011010110101101101011010010000100001000010000100001000110111101101000010000100001000010000100011011110111011111011110110100001000010000100001000010000100001000010000100001000110101001110011101101100111001011000110001100"),
                ("1100111001100111011010110100111011010110101101101011010010000100001000010000100001000110111101101000010000100001000010000100011011110111011111011110110100001000010000100001000010000100001000010000100001000110101001110011101101100111001011000110001100"),
                ("1100111001110011100111001110011001110011101101101011010010000100001000010000100001000010000100001000010000100010111110111101110111101111011110111101110100001001010010100001000010000100001000010000100101001100111001110011110010110001100011001100111001"),
                ("1101011010011001100111001110011011010110100111101011010010010100101000010000100001000010000100011011101111011100001000010000100001000011101100001000010100001001010010100101000010000100001000010000100101001100111001110011100111111011110011001111111111"),
                ("1101011010011001100111001110011011010110100111101011010010010100101000010000100001000010000100011011101111011100001000010000100001000011101100001000010100001001010010100101000010000100001000010000100101001100111001110011100111111011110011001111111111"),
                ("1111111111111111100111001110011011010110101100100101001010000100001000010000100001000110111101100001000010000100001000010000111011110111101100001000011101101000010000100001001010010100101001010010100001000110101001110011100111001110011111111111111111"),
                ("1111111111111111100111001100111001110011100110100001000010000100001000010000100001000010000100001000101111011110111110111101111011110111011100001000011011101000010000100001000010000100111000110001101011010110001001110011100111100111001111111111111111"),
                ("1111111111111111100111001100111001110011100110100001000010000100001000010000100001000010000100001000101111011110111110111101111011110111011100001000011011101000010000100001000010000100111000110001101011010110001001110011100111100111001111111111111111"),
                ("1111111111111111101011010110000100101001010000100001000010010100101000010000100001000010000100001000110111101111011101111011100001000010000100001000011011101000010000100101001010011100001001010010100101001110001001110011100111100111001011001111111111"),
                ("1111111111111110100101001010010100101001010000100001000010000100001000010000100001000101111011110111101111011110111000010000100001000010000110111101111101101000010000100101001010011100011000110000100101001100111100111001110011100111001110011100111001"),
                ("1111111111111110100101001010010100101001010000100001000010000100001000010000100001000101111011110111101111011110111000010000100001000010000110111101111101101000010000100101001010011100011000110000100101001100111100111001110011100111001110011100111001"),
                ("1111111111111111001110011100111001110011110100100001000010000100001000010000100001000110111101100001000010000110111000010000110111101111011111011110111101101000010000100001000010000100101001010011101011010100111011010110100111100111001110011100111001"),
                ("1111111111111111011010110101101011010110100111100011000010010100101000010000100001000110111101100001000010000100001000010000111011110110100010111101111011101000010000100001000010000100001000010000100101001101101011010110100111100111001110010110001100"),
                ("1111111111111111011010110101101011010110100111100011000010010100101000010000100001000110111101100001000010000100001000010000111011110110100010111101111011101000010000100001000010000100001000010000100101001101101011010110100111100111001110010110001100"),
                ("0001100011011001011010110101101011010110101101001110011010010100101000010000100001000101111011100001000010000100001000010000100001000010000111011110110000111011110110100001000010000100001000010000100001000100111011010110101100110001100111101111011110"),
                ("0001100011011001011010110101101011010110101101001110011010010100101000010000100001000101111011100001000010000100001000010000100001000010000111011110110000111011110110100001000010000100001000010000100001000100111011010110101100110001100111101111011110"),
                ("1101011010111011011010110101101001110011101101101011010010010100101000010000100001000010000100010111000010000100001000010000100001000010000111011110110000111011110110100001000010000100001000010000100101001101101001110011101101111011110111100110001100"),
                ("1100111001110011011010110100111001110011100111100011000010000100001000110111101110111101111011100001000010000100001000010000100001000010000110111101111011101000010000100001000010000100001000010000100001000100111001110011100110110001100111111111111111"),
                ("1100111001110011011010110100111001110011100111100011000010000100001000110111101110111101111011100001000010000100001000010000100001000010000110111101111011101000010000100001000010000100001000010000100001000100111001110011100110110001100111111111111111"),
                ("1100111001110011001110011101101011010110110000100101001010000100001000110111101100001000010000100001110111101110111000010000100001000010000100001000010000110111101110100001000010000100001000010000100001000110001001110011110011110111101111111111111111"),
                ("1111011110111011100111001101101001110011010010100001000010010100101000010000100011011000010000100001101111011100001110111101100001000010000100001000010000110111101111011101000010000100001001010010100101001100111001110011011000111001110111111111111111"),
                ("1111011110111011100111001101101001110011010010100001000010010100101000010000100011011000010000100001101111011100001110111101100001000010000100001000010000110111101111011101000010000100001001010010100101001100111001110011011000111001110111111111111111"),
                ("1111111111011100110001100110011001110011010011101011010010010100101000010000100001000101111011100001101111011110111110111101101000010000000110111101110100001000010000100001000010000100001001010011100011000110101001110011110011100111001111111111111111"),
                ("1111111111111110110001100111010110001100110101001110011010010100101000010000100001000101111011111011010000100011011110111101101000010001011110111101110100001000010000100001000010000100001001010011100011000010011100011000100111011010110111111111111111"),
                ("1111111111111110110001100111010110001100110101001110011010010100101000010000100001000101111011111011010000100011011110111101101000010001011110111101110100001000010000100001000010000100001001010011100011000010011100011000100111011010110111111111111111"),

                -- 6_explosion_3_1
                ("1111111111111111111011110110011100111001110100001100011111111111111111111111111111111111111111111111110101101011001110011100101100011001011011001110011101011001110011100101100011001111111111111111111111111111111111111111111111110111101011001011010110"),
                ("1111111111111111111011110110011100111001110100001100011111111111111111111111111111111111111111111111110101101011001110011100101100011001011011001110011101011001110011100101100011001111111111111111111111111111111111111111111111110111101011001011010110"),
                ("1111111111011101110111101110011100111001111010110001100111111111111111111111111111111111111111111111011000110011001100111001110011100111100111001110011100111001110011001110110101101111111111111111111111111111111111111111111111111011110110011001110011"),
                ("0110001100011001100111001100111011010110101101011010110101101011010011010010100111010110011100111001110011100111001101101011011001110011100110110101101011010110101101001110011100111011010011100110110001100110011110111101011000110001100110011001110011"),
                ("0110001100011001100111001100111011010110101101011010110101101011010011010010100111010110011100111001110011100111001101101011011001110011100110110101101011010110101101001110011100111011010011100110110001100110011110111101011000110001100110011001110011"),
                ("1110111101110011011010110101101001110011101101011010110101101011010011010010100111000100111001111001110011100111001100111001110110101101011010011100111101010011100111101011010110101011010110101101011010110101101100111001110011001110011100111011010110"),
                ("0110001100100111001110011101101001110011100111011010110101101011010011010010100101001100111001110110101101011010011101101011010110101101011011010110100100101001010010100110011100111011010110101101011010110110011100111001110011011010110100111011010110"),
                ("0110001100100111001110011101101001110011100111011010110101101011010011010010100101001100111001110110101101011010011101101011010110101101011011010110100100101001010010100110011100111011010110101101011010110110011100111001110011011010110100111011010110"),
                ("1101011010010010100101001110001001110011101101011010110100111001111010010000100001000100111001110110100111001110110101101011010011100111011010011100111100001001010010100111010110101001110011100111001110011110101101011010100111001110011101101011010110"),
                ("1001110011110100100001000010011100011000110101001110011110001100001000010000100001000010000100001001110101101011010110101101011000110001101011000110000100001000010000100111000110000100101001010010100001000010000100101001010010100101001100111011010110"),
                ("1001110011110100100001000010011100011000110101001110011110001100001000010000100001000010000100001001110101101011010110101101011000110001101011000110000100001000010000100111000110000100101001010010100001000010000100101001010010100101001100111011010110"),
                ("0100101001010010100101001010000100001000010010100101001010010100101000010000100001001010000100001000010010100101000010000100001001010010100001001010010100001000010000100001001010010100111000110000100101001010010100101001010000100001000100111011010110"),
                ("0100101001010010100101001010000100001000010010100101001010010100101000010000100001001010000100001000010010100101000010000100001001010010100001001010010100001000010000100001001010010100111000110000100101001010010100101001010000100001000100111011010110"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001010010100101000010000100001001010011100001001010010100001000010010100001000010000100001000100111011010110"),
                ("0100001000010000100001000110111101111011010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100001000010000100001000010000100001001010010100101001010010100101001010010100001000010000100001000110101001110011"),
                ("0100001000010000100001000110111101111011010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100001000010000100001000010000100001001010010100101001010010100101001010010100001000010000100001000110101001110011"),
                ("0100001000010001101111011000011011110111010000100001000010000100001000010000100001000010000100001000010000100001000010000100011011110110100001000010000100001000010000100001000010000100001000010000100101001010010100001000010000100001000010010100101001"),
                ("1011110111101110000100001000011011110111010001011110111110111101111011101111011101000010000100011011010000100001000110111101110111101110100011011110111101101000010000100001000010000100001000010000100101001010000100001000101011101111011010000100001000"),
                ("1011110111101110000100001000011011110111010001011110111110111101111011101111011101000010000100011011010000100001000110111101110111101110100011011110111101101000010000100001000010000100001000010000100101001010000100001000101011101111011010000100001000"),
                ("1101111011000010000100001000010000100001101110000100001000010000100001101111011101000010000100000001110111101101000010000100011011110111101100001000010000110111101111011111011110110100001000010001101111011010000100001000101110000100001110110100001000"),
                ("0100001000101111011110111110110000100001000010000100001000010000100001101111011111011101111011100001101111011101000010000100010111101110000100001000010000100001000010000110111101111101100001000011011110111101111011110111000010000100001101110100001000"),
                ("0100001000101111011110111110110000100001000010000100001000010000100001101111011111011101111011100001101111011101000010000100010111101110000100001000010000100001000010000110111101111101100001000011011110111101111011110111000010000100001101110100001000"),
                ("1101111011101110000100001101110000100001000010000100001000010000110111101111011111011101111011100001000010000110111010000100001000010001011100001000010000100001000010000100001000010000110111101110000100001000011101111011101110000100001000010100001000"),
                ("1101111011110111101111011000010000100001000010000100001000010000100001000010000110111110111101100001000010000111011010000100001000010001011100001000010000100001000010000100001000010000111011110111101111011000010000100001101111101111011110110100001000"),
                ("1101111011110111101111011000010000100001000010000100001000010000100001000010000110111110111101100001000010000111011010000100001000010001011100001000010000100001000010000100001000010000111011110111101111011000010000100001101111101111011110110100001000"),
                ("0100001000010000000100001000010000100001000010000100001110111101110111000010000100001110111101111011000010000110111110111101101000010001011110111101111011100001000011101110111101111011100001000011011110111000010000100001101110100001000010000100001000"),
                ("0100001000010000000100001000010000100001000010000100001110111101110111000010000100001110111101111011000010000110111110111101101000010001011110111101111011100001000011101110111101111011100001000011011110111000010000100001101110100001000010000100001000"),
                ("1011110111000010000100001000010000100001000010000100001010000100010111000010000100001101111011111011110111101110111101111011111011110111011100001000010000100001000010100011011110110000100001000011011110111101110000100001000011011110111010000100001000"),
                ("1011110111101110000100001000011011110111110111101111011101111011111011101111011100001000010000100001000010000110111110111101110111101111011101000010001011100001000011011100001000010000100001000010000100001000010000100001000010000100001110110100001000"),
                ("1011110111101110000100001000011011110111110111101111011101111011111011101111011100001000010000100001000010000110111110111101110111101111011101000010001011100001000011011100001000010000100001000010000100001000010000100001000010000100001110110100001000"),
                ("0100001000010000000100001000011011110111000010000100001101111011111011110111101110111101111011111011010000100001000010000100011011110110100011011110110000110111101110000110111101111011110111101110000100001000010000100001101111011110111110110100001000"),
                ("0100001000010001011110111101110100001000110111101111011010000100001000010000100001000010000100001000010010100101001010000100001000010000100011011110111101101000010000000101000010000100010111101110000100001000011011110111110110100001000010000100101001"),
                ("0100001000010001011110111101110100001000110111101111011010000100001000010000100001000010000100001000010010100101001010000100001000010000100011011110111101101000010000000101000010000100010111101110000100001000011011110111110110100001000010000100101001"),
                ("0100001000010001011110111010000100001000010000100001000010000100001000010010100101001010000100001000010010100101000010000100001000010000100001000010000100001000010001011111011110110100001000010001011110111110110100001000010010100001000010000100101001"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010010100101001010000100001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010100001000010001101011010"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010010100101001010000100001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010100001000010001101011010"),
                ("0100001000010000100001000010000100001000010000100001000010000100001001110001100011000010010100101001010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010010100101001010010100101001010000100001000"),
                ("0100101001010010100101001010000100001000010000100001000010000100001001110001100001001110001100001001010000100001000010000100001001010010100101001010010100101000010000100001000010000100001001010010100101001010010100001000010000100001000010000100001000"),
                ("0100101001010010100101001010000100001000010000100001000010000100001001110001100001001110001100001001010000100001000010000100001001010010100101001010010100101000010000100001000010000100001001010010100101001010010100001000010000100001000010000100001000"),
                ("1100011000110000100101001010000100001000010010100001000010010100111010010010100101001110101101001000010010100101001010000100001001010010100111000110000100101001010010100001001010011101001001010011100011000110001100011000110000100101001010000100001000"),
                ("1100011000110000100101001010000100001000010010100001000010010100111010010010100101001110101101001000010010100101001010000100001001010010100111000110000100101001010010100001001010011101001001010011100011000110001100011000110000100101001010000100001000"),
                ("0100101001110101001110011110001001110011101101001110011101101011010011100111001111000110001100011010100111001110011110101101011010110101101010011100111101011010110100100110011100111011010011100111001110011101101001110011110100100101001010000100101001"),
                ("1100011000100111001110011100111001110011100111011010110101101011010110110011100110011100111001110011100111001110011100111001111010110101101010110101101011010110101101101010011100111011010110101101011010110110011011010110110100100101001010011001110011"),
                ("1100011000100111001110011100111001110011100111011010110101101011010110110011100110011100111001110011100111001110011100111001111010110101101010110101101011010110101101101010011100111011010110101101011010110110011011010110110100100101001010011001110011"),
                ("1001110011110010110001100110011001110011101101011010110100111001110011110011100110011100111001110011100111001111001101101011010011100111001110110101101011010110101101100110011100111011010110101101001110011110011001110011100111101011010010011001110011"),
                ("1011010110110010111001110111010110001100111100110001100110011100111001110011100111001110011100110011111101111001100110011100110011100111011010110101101011010110101101100111001110011011011001110011100111001110011100111001110011100111001100111100111001"),
                ("1011010110110010111001110111010110001100111100110001100110011100111001110011100111001110011100110011111101111001100110011100110011100111011010110101101011010110101101100111001110011011011001110011100111001110011100111001110011100111001100111100111001"),
                ("1111111111111111111111111111111111111111111101111011110110011100111001110011100101100111111111111111011000110001100011000110011001110011111111111111111111111111111111100111001110011001101100011001111011110011001111111111111111100111001110010110001100"),
                ("1111111111111111111111111111111111111111011001111011110011000110011001110011100111111111111111111111111111111111001011000110011101111011111111111111111111111111111111111111001110011100101100011000111001110111111111111111111111111111111110010110001100"),
                ("1111111111111111111111111111111111111111011001111011110011000110011001110011100111111111111111111111111111111111001011000110011101111011111111111111111111111111111111111111001110011100101100011000111001110111111111111111111111111111111110010110001100"),

                -- 7_explosion_0_0
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000110011001011000110011001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000110011001011000110011001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110010110011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110010110011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111110011100111001110011100110011110011100111001110011100111001110011100111001110011100110011100111001111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110110011100111001110011100110110110011100111001110011100111001110011100111001110011100110011100111001110110101101001111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110110011100111001110011100110110110011100111001110011100111001110011100111001110011100110011100111001110110101101001111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110110001100110011100111001100111001111001110011100111001110011100111001110011100111001110011011010110101101011010110101101001111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110110001100110011100111001100111001111001110011100111001110011100111001110011100111001110011011010110101101011010110101101001111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001110011100110011100111001111001100111001111001110011100110011110011100111001110011011010011100111001110011100111100111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001110011100110110110011100111001110011100110011100111001110011100111100110011100111100110011100111001111001110011100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001110011100110110110011100111001110011100110011100111001110011100111100110011100111100110011100111001111001110011100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100011001100111001110011100111001110011100110011100111001111001110011100110110101101011010110101101011010110101101100110011100111001110110101101011011001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001110011100110011100111001110110110011100110110101101011010110101101011010110101101011010110101101011010110101101001111001110011100111001110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001110011100110011100111001110110110011100110110101101011010110101101011010110101101011010110101101011010110101101001111001110011100111001110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001110011100111001100111001110110100111001111010100111001110110101101001110011100111011010110101101011010110101101001111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110011110011100110011110101101010110110101101001001010010100111000110000100110011100111011010110101101011010011100111100111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100110011110011100110011110101101010110110101101001001010010100111000110000100110011100111011010110101101011010011100111100111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001100111001110110100111001110110110101101001001110001100001001010010100111010110101001110110101101001111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001110011100110011101101011010011110001100001001010010100101001010011101001001010010100111010110101001111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001110011100110011101101011010011110001100001001010010100101001010011101001001010010100111010110101001111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100111001101101011010011110001100001001010010100101001010011101010011100111101011010110101001110011100111001111001110011100111001110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100111001101101011010011110001100001001010010100101001010011101010011100111101011010110101001110011100111001111001110011100111001110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001101101011010011110011100110110101101011010011010010100101001110101101010011100111011010110101101011010110101101001110011100111011010110101101011010110110011110111101111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011001110011101101011010110110011100110110101101011011010010010100101001110101101010011100111101010011100111011010011100111101010011100111011010011100111001110011110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011001110011101101011010110110011100110110101101011011010010010100101001110101101010011100111101010011100111011010011100111101010011100111011010011100111001110011110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011001110011101101011010110101101011010110101101011010011110101101001001100111001111010110101100011010110101001110011100111011010011100111100111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001101101011010110101101011010110101101011011010110101101011010100111001111010110101001111010110100100110011100111011011001110011100111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001101101011010110101101011010110101101011011010110101101011010100111001111010110101001111010110100100110011100111011011001110011100111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100110110101101011010110101101011010011110001100010011100111001111010110101001110011100111001110110101101011010011100111100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111101100111001110011100111001101101011010110101101011010110100111001110011110001100001001010010100110011100111001110011100111011010110101101100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111101100111001110011100111001101101011010110101101011010110100111001110011110001100001001010010100110011100111001110011100111011010110101101100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011101111011110011000110011001110011100110011101101011010110101101011011000010010100101001010011100010011100111001110011100111011010110101101100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111101111011110111101111011001110011100110011101101011010110100111001101001010010100101001010011100010011100111101010011100111001110011100111011010011100111100111001111011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111101111011110111101111011001110011100110011101101011010110100111001101001010010100101001010011100010011100111101010011100111001110011100111011010011100111100111001111011111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111101100111001110011100111001100111001110011101101011010011110001100001001010010100111010110101101011010110101001110011100111001110011100111011010110101101100111001111101111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111101100111001110011100111001100111001110011101101011010011110001100001001010010100111010110101101011010110101001110011100111001110011100111011010110101101100111001111101111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110011001100111001110011100110011101101011010011101101011010110110101101001001110001100011010110101100011000110001101010011100111001110011100111001111001110011100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001100111001110011100110011101101011010110100111001110011100111001111010110001100011010110101101011010110101101011010110101101010011100111001110011100111100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001100111001110011100110011101101011010110100111001110011100111001111010110001100011010110101101011010110101101011010110101101010011100111001110011100111100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011000110001100110011100110011101101011010011110101101010011101101011011010010010100111010110101101011000110001100011010110101101010011100111001110011100110110001100111101110111101111111111111111111111111111111"),
                ("1111111111111111111111111111101111011110111101100111001110011100111001101101011010110100111001110110100111001111000010010100101001010011101010011100111101011010110101100011010110101001110011100111100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111101111011110111101100111001110011100111001101101011010110100111001110110100111001111000010010100101001010011101010011100111101011010110101100011010110101001110011100111100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001100111001110011100110011100111001110011100111001110110100111001111010010010100111000110001101011010110101101010011100111101011010110101001110011100111100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001100111001110011100111001011000110010011100111001110011100111001111010110101101011000110001101011010110101001110011100111001110011100111001111001110011111011110111101110111101111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001100111001110011100111001011000110010011100111001110011100111001111010110101101011000110001101011010110101001110011100111001110011100111001111001110011111011110111101110111101111111111111111111111111111111"),

                -- 7_explosion_0_1
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0111001110011101111011110011100111001110111101111011110111101111011111111111111101100110011100111001110011100111111111111111111001110011100111001110010110011001110010110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0111001110011101111011110011100111001110111101111011110111101111011111111111111101100110011100111001110011100111111111111111111001110011100111001110010110011001110010110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0110001100011001111011110011000110001100011001111011110111101111001110111101111011001110011100111001110011100111001110011100111001110011100111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001011001100111001110011100111001111101111011110110011100111001110011100110011100111001111001110011100111001110011100111001110011100111001110011100111001110011100101100011001111011110111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001011001100111001110011100111001111101111011110110011100111001110011100110011100111001111001110011100111001110011100111001110011100111001110011100111001110011100101100011001111011110111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001110011100111001110011100111001111101111001100110011100111001101101011010110101101011010110110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1100111001110011100111001110011100111001110011100111001111101111001100110011100111001101101011010110101101011010110110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1100111001100111100111001100111001110011100111100111001110011100111001110011100110110101101011010110101101011010011110011100111001110011100110011100111100111001110011100111001110011001111001110011100111001110011100111001111111111111111111111111111111"),
                ("0110001100100111011010110101101011010110101101001110011110011100111001101101011010110101101011010110110011100111001110011100111001110011001111001110011100111001110011100111001110011001110011100111100111001110011100111001111111111111111111111111111111"),
                ("0110001100100111011010110101101011010110101101001110011110011100111001101101011010110101101011010110110011100111001110011100111001110011001111001110011100111001110011100111001110011001110011100111100111001110011100111001111111111111111111111111111111"),
                ("1001110011100111011010110100111011010110100111001110011100111001110011101101011010110101101011010110101101011010110110011100110011100111011010011100111100110011100111001110110101101100111001110011011010110100111100111001111111111111111111111111111111"),
                ("1001110011100111001110011110101001110011101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101001111010110101001110011100111001111001110011001111001110011100111001110011100111001110011111111111111111111111111"),
                ("1001110011100111001110011110101001110011101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101001111010110101001110011100111001111001110011001111001110011100111001110011100111001110011111111111111111111111111"),
                ("1001110011101101011010110100111001110011101101001110011101101011010110101101011010011110101101010011110101101010011100111001110011100111011010110101101011010110101101100111001110011100111001110011100111001110011100111001110011111011110111111111111111"),
                ("1001110011100111001110011101101001110011110101100011000100111001110110100111001111000110101101011010010010100101001110001100011000110001101011010110101001111001110011100111001110011100111001110011100111001110011100111001110010110001100111111111111111"),
                ("1001110011100111001110011101101001110011110101100011000100111001110110100111001111000110101101011010010010100101001110001100011000110001101011010110101001111001110011100111001110011100111001110011100111001110011100111001110010110001100111111111111111"),
                ("1101011010110101100011000110101101011010010010100101001010010100111000100111001110011110101101001001010010100101001010010100101001010010100101001010011101010110101101011010011100111001111001110011100111001110011100111001110011100111001111111111111111"),
                ("1101011010010010100101001010011100011000110000100101001010010100101001110001100010011100111001110011110101101011010010010100101001010011100001001010011001110110101101011010011100111100111001110011100111001110011100111001110010110001100111111111111111"),
                ("1101011010010010100101001010011100011000110000100101001010010100101001110001100010011100111001110011110101101011010010010100101001010011100001001010011001110110101101011010011100111100111001110011100111001110011100111001110010110001100111111111111111"),
                ("1100011000110000100101001110101101011010110101101011010010010100101001010010100111010110101101011010100111001110011010010100101001010010100111000110001011010110101101011010011100111100111001110011100111001110011100111001110011100111001111111111111111"),
                ("1100011000110000100101001110101101011010110101101011010010010100101001010010100111010110101101011010100111001110011010010100101001010010100111000110001011010110101101011010011100111100111001110011100111001110011100111001110011100111001111111111111111"),
                ("1101011010110101101011010110101101011010110001101011010110001100011000010010100110011100111001111000110101101010110110101101011010110100100101001010011001110110101101011011001110011011010110101101100111001110011100111001110011100111001111111111111111"),
                ("1101011010110101001110011110001101011010110001101011010100111001110011100111001110011110101101011010100111001110110100111001101001010011101010011100111001110110101101011010011100111001110110101101001110011100111100111001110011100111001111111111111111"),
                ("1101011010110101001110011110001101011010110001101011010100111001110011100111001110011110101101011010100111001110110100111001101001010011101010011100111001110110101101011010011100111001110110101101001110011100111100111001110011100111001111111111111111"),
                ("1001110011110101101011010110001101011010110101001110011110101101010011100111001110011010010100110011101101011010110110101101001001010011001110110101101011010110101101100111001110011001110110101101001110011100111100111001110011100111001111111111111111"),
                ("1001110011100111101011010110101101011010100111001110011100111001110011100111001110110100111001110011100111001110110110101101011010110101011010110101101011010110101101001110011100111001110110101101011010110110011100111001110011111111111111111111111111"),
                ("1001110011100111101011010110101101011010100111001110011100111001110011100111001110110100111001110011100111001110110110101101011010110101011010110101101011010110101101001110011100111001110110101101011010110110011100111001110011111111111111111111111111"),
                ("1001110011110101100011000110101101011010100111001110011100111001110110101101011010110101101011010110110101101010011100111001110011100111001110110101101011010110101101001110011100111100110011100111001110011110011100111001111111111111111111111111111111"),
                ("1001110011110101101011010100111001110011100111001110011100111001110110101101011010011110011100110011100111001110011100111001111001110011100110011100111011010110101101011011001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1001110011110101101011010100111001110011100111001110011100111001110110101101011010011110011100110011100111001110011100111001111001110011100110011100111011010110101101011011001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1001110011100111001110011100111001110011100111011010110101101011011001110011100111001110011100111001101101011010110100111001111001110011100111001110011001110011100111011011001110011100111001110011100111001011000110001100111111111111111111111111111111"),
                ("1100111001100111001110011100111001110011110011011010110100111001111001110011100111001110011100111001100111001110110110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1100111001100111001110011100111001110011110011011010110100111001111001110011100111001110011100111001100111001110110110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111011110110011100111001011001100111001110011100111001110011100111001110011100111001110011100111001100111001110110110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111011110110011100111001011001100111001110011100111001110011100111001110011100111001110011100111001100111001110110110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111011110110010110001100111101100111001011001111011110111011110101100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110010110001100011001111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1110111101110010110001100111011100111001011001111011110111101111011111111111111111001011000110001100011000110011101111011110111111111111111101100011000110011101111010111011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1110111101110010110001100111011100111001011001111011110111101111011111111111111111001011000110001100011000110011101111011110111111111111111101100011000110011101111010111011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_0_2
                ("1111111111111111111111111111111110111101111101111011110110011100110011100111001110011100111001110011110101101011010110001100011010110101101010011100111001110011100111001101100011001100111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101111101111011110110011100110011100111001110011100111001110011110101101011010110001100011010110101101010011100111001110011100111001101100011001100111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001100111001110011110101101011010100111001111010110101101011010110001100001001010011101010011100111011010011100111001110011100111001111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100011001100111001100111001110011110101101011000110101101011010100111001111010010010100101001010011100010011100111011010011100111011010110101101100111001110011100111001111101111011110111101111111111111111111111111"),
                ("1111111111111111111111111111110110001100011001100111001100111001110011110101101011000110101101011010100111001111010010010100101001010011100010011100111011010011100111011010110101101100111001110011100111001111101111011110111101111111111111111111111111"),
                ("1111111111111111111111111111111110111101111100110001100100111001110011100111001111010110101101011000110001100011010110101101001001010011101010110101101001111010110101001110110101101001111001110010110001100011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001100111001110011100111001111010110101101011010110101101011010110101101011000110001101010011100111001110011100111011010110101101001111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001100111001110011100111001111010110101101011010110101101011010110101101011000110001101010011100111001110011100111011010110101101001111001110011100111001011000111001110111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100011001100111001110011100110011100111001110011100111001111010110001100011000110101101011000110000100111010110101011010110101101001110110101101001111001110011100111001011001111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111101100111001101101011010110100111001110011100111001110011110101101011010110101101001001010010100111000110001001110110101101001110011100111100111001110011100111001111101111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111101100111001101101011010110100111001110011100111001110011110101101011010110101101001001010010100111000110001001110110101101001110011100111100111001110011100111001111101111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111011100111001100111001110110100111001110011100111001111010100111001111000010010100101001010010100110011100111011010110101101001111001110011100111110111101111011110111101111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111011110111011100111001100111001110110100111001110011100111001111010100111001111000010010100101001010010100110011100111011010110101101001111001110011100111110111101111011110111101111011110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001101101011010110100111001110011100111001111000010010100101001010011100010110101101011010110101101001111001110011100101100011001111011110011101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001101101011010110100111001110011100111001101001010010100111000110001001110011100111011010110101101011010110101101100111001110011100111001111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001101101011010110100111001110011100111001101001010010100111000110001001110011100111011010110101101011010110101101100111001110011100111001111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001100111001110110101101011010011100111001110011110101101010011100111001111000110001001110110101101011010110101101011011001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001110011100110110100111001101001110101101010011110101101010011100111101011010110101101010110101101011010110101101011010110101101100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001110011100110110100111001101001110101101010011110101101010011100111101011010110101101010110101101011010110101101011010110101101100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001100111001110110100111001110011110101101011000110101101010011100110100111010110101001110110101101011010110101101011010110101101001110011110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011001110011100111001110110100111001111010100111001110110100111001111010100111001111010110100100101001010011101010110101101011011001110011011010110101101001110011110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011001110011100111001110110100111001111010100111001110110100111001111010100111001111010110100100101001010011101010110101101011011001110011011010110101101001110011110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101110011011010110101101011010110100111001110011101101011010110101101011010110100111001111010110100100101001010011001110110101101011011001110011001110110101101100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101110011100111001110011100110011100111001110011110101101011010100111001111010010010100101001010010100111000110001001110110101101100111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101110011100111001110011100110011100111001110011110101101011010100111001111010010010100101001010010100111000110001001110110101101100111001110011100111001110011100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100110011110101101001001010010100111010010010100101001010010100111000110001001110110101101001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100110011110101101001001010010100111010010010100101001010010100111000110001001110110101101001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100110011101101011010011110101101001001010010100111000110000100111010110101011010011100111011010011100111100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001100111001110110101101011010110100111001101001110001100001001010010100111010110101011011010110101001111001110011001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100111001100111001110110101101011010110100111001101001110001100001001010010100111010110101011011010110101001111001110011001111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011100111001110011100110011101101011010110101101011010110100111001110011101101011010011100111101010011100111011010011100111100111001110011100111001110011100111001110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101110011100111001110011100110011101101011010110101101011010110101101011010110101101011010110101101011011001110011011010011100111001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111111110111101110011100111001110011100110011101101011010110101101011010110101101011010110101101011010110101101011011001110011011010011100111001111001110011100111001110011100111001110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110011001100111001110011100110110101101011010011100111001111001101101011010110101101011010110101101011011001110011100110011100111001111001110011100111001110011100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001110011100110011100111001111001100111001111001100111001110011100111001111001110011100111001110011011011001110011100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001110011100110011100111001111001100111001111001100111001110011100111001111001110011100111001110011011011001110011100111001110011100111001011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100111001100111001110011100111001110110110011100111001110011001111001110011100110011100111100110011100111001111001110011100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100110011101101011010110101101011010110110011100111001110011100111001110011100111001110011100110011100111100111001110010110001100111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100110011101101011010110101101011010110110011100111001110011100111001110011100111001110011100110011100111100111001110010110001100111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100110011101101011010011100111001111001110011100111001110011100111001110011100111001110011011011001110011100111001110011111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100110011101101011010011100111001111001110011100111001110011100111001110011100111001110011011011001110011100111001110011111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111011000110001100110011100111001110011100110011100111001111001110011100111001110011100111001110011100111001110011001111001110011100111001110011111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111101100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111101100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100101100011001100101100011001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100101100011001100101100011001111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_0_3
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011110101100011000110011111111111111111101111011110101100011000110001100011001100111111111111111111110111101111011110011001100111001111010110001100110011110111101"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011110101100011000110011111111111111111101111011110101100011000110001100011001100111111111111111111110111101111011110011001100111001111010110001100110011110111101"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111011000110001100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110010110011101111011111011110011001100111001111100110001100110011111011110"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011011010011100111100111001110011100111001110011100111001110011100111001110011100111001011001100111001110011111011110"),
                ("1111111111111111111111111111111111111111111111100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011011010011100111100111001110011100111001110011100111001110011100111001110011100111001011001100111001110011111011110"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011011010011100111100111001110011100111001110011100110011100111011010110110011001110011100111001110011100111100111001"),
                ("1111111111111111111111111111111111111111011001100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011011010011100111100111001110011100111001110011100110011100111011010110110011001110011100111001110011100111100111001"),
                ("1111111111111111111111111111110110001100011001100111001110011100111001110011100110110100111001110011110011100111001110011100110011100111011010110101101100111001110011100111001110011100110110101101011010110100111001110011100111001110011100111001110011"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001110011100110110101101011010110100111001111001110011100110011100111001110011100111001111001110011001110110101101011010011100111001110011100111001110011100111101011010110101001110011"),
                ("1111111111111111111111111111111100111001110011100111001110011100111001110011100110110101101011010110100111001111001110011100110011100111001110011100111001111001110011001110110101101011010011100111001110011100111001110011100111101011010110101001110011"),
                ("1111111111111111111111111111111100111001110011001110011100111001111001100111001110011101101011010110101101011010011100111001110011100111001111010110101011010110101101011010110101101011010011100111001110011100111101011010110101100011000110101001110011"),
                ("1111111111111111111111111110011100111001110011011010110101101011010011100111001110011101101011010110101101011010110110101101011010110101011010011100111001110011100111011010011100111001110011100111001110011100111101011010110101101011010100111001110011"),
                ("1111111111111111111111111110011100111001110011011010110101101011010011100111001110011101101011010110101101011010110110101101011010110101011010011100111001110011100111011010011100111001110011100111001110011100111101011010110101101011010100111001110011"),
                ("1111111111111111100111001110011100111001100111001110011101101011010011110011100111001101101011010110101101011010011010010100111010110101011010110101101001101001010011001110011100111001111010110101001110011110101101011010110001101011010110101001110011"),
                ("1111111111111111100111001110011100111001100111001110011101101011010011100111001110110101101011010011100111001111010010010100110011100111011010011100111101011010110101001110011100111001110011100111101011010110001101011010110001001110011110101101011010"),
                ("1111111111111111100111001110011100111001100111001110011101101011010011100111001110110101101011010011100111001111010010010100110011100111011010011100111101011010110101001110011100111001110011100111101011010110001101011010110001001110011110101101011010"),
                ("1111111111111111100111001110011100111001110011100111001101101011010110110011100110110101101011010011010010100101001110101101011010110101011011010110101100010011100111001101001010011100011000110001101011010110001101011010110101101011010110101101011010"),
                ("1111111111111111100111001110011100111001110011100111001110011100111001100111001110110101101011010110110001100001001010010100101001010011001110011100111101011010110101101001001010010100101001010011101011010110101101011010110100100101001110001100011000"),
                ("1111111111111111100111001110011100111001110011100111001110011100111001100111001110110101101011010110110001100001001010010100101001010011001110011100111101011010110101101001001010010100101001010011101011010110101101011010110100100101001110001100011000"),
                ("1111111111111110110001100110011100111001110011100111001110011100111001100111001110110101101011010011010010100111000010010100101001010011101011010110101001110011100111001111000110000100101001010010100101001110001100011000010010100101001010011101011010"),
                ("1111111111111110110001100110011100111001110011100111001110011100111001100111001110110101101011010011010010100111000010010100101001010011101011010110101001110011100111001111000110000100101001010010100101001110001100011000010010100101001010011101011010"),
                ("1111111111111111100111001110011100111001110011100111001110011100110011100111001110110101101011011010010010100101001010010100101001010010100101001010010100111010110101001110011100111100001001010010100101001010011101011010110101100011000110101101011010"),
                ("1111111111111110110001100110011100111001110011100111001110011100111001110011100111001110011100110011110101101011010110001100011000110000100101001010011101011010110101100010011100111011010011100111100011000110101001110011101101001110011100111001110011"),
                ("1111111111111110110001100110011100111001110011100111001110011100111001110011100111001110011100110011110101101011010110001100011000110000100101001010011101011010110101100010011100111011010011100111100011000110101001110011101101001110011100111001110011"),
                ("1111111111111111111011110110011100111001110011100111001110011100111001110011100111001101101011010110101101011010110100111001110011100111001111010110101001111010110101001110110101101011010110101101001110011101101001110011100111011010110101101001110011"),
                ("1111111111111111111111111110011100111001110011100111001110011100110011110011100110011100111001110011110101101010011101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101001110011110101001110011100111001110011"),
                ("1111111111111111111111111110011100111001110011100111001110011100110011110011100110011100111001110011110101101010011101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101001110011110101001110011100111001110011"),
                ("1111111111111111111111111111111100111001100111011010110110011100111001101101011010011100111001111001100111001110110100111001111001110011011010110101101011010110101101011010110101101001110011100111001110011100111011010110100111011010110100111001110011"),
                ("1111111111111111111111111111111100111001110011100111001100111001110011110011100111001110011100111001110011100110011110011100111001110011100111001110011011010110101101011010110101101100111001110011001110011101101011010110101101011010110100110110001100"),
                ("1111111111111111111111111111111100111001110011100111001100111001110011110011100111001110011100111001110011100110011110011100111001110011100111001110011011010110101101011010110101101100111001110011001110011101101011010110101101011010110100110110001100"),
                ("1111111111111111111111111111111100111001110011100111001110011100110011110011100111001110011100111001100111001111001110011100111001110011001110110101101011010110101101011011001110011100111001110011100111001100111001110011100111100111001100111100111001"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011011010110101101011010110101101100111001110010110011110111101100111001110011100111001110011100111001110011100111001"),
                ("1111111111111111111111111111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011011010110101101011010110101101100111001110010110011110111101100111001110011100111001110011100111001110011100111001"),
                ("1111111111111111111111111111111111111111111111111011110011000110011001110011100111001110011100111001110011100111001110011100111001110011100110011100111001111001110011100111001110011111011110111101100111001110011100111001011001100111001110011100111001"),
                ("1111111111111111111111111111111111111111111111111011110011000110011001110011100111001110011100111001110011100111001110011100111001110011100110011100111001111001110011100111001110011111011110111101100111001110011100111001011001100111001110011100111001"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111011000110001100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111110111100111011110111101111011110011000110001100011001111011110011000110001100"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111101100110011100101100110011100111001110011100111111111111111111001110011100111001110010110011111111111111111110111101111011110111100111001110011101111011110011100111001110"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111101100110011100101100110011100111001110011100111111111111111111001110011100111001110010110011111111111111111110111101111011110111100111001110011101111011110011100111001110"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_1_0
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010110101001111010110101001110011100111001111001110011111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011010110101001111010110101001110011100111001111001110011111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100111001110011110011100101100011000110011110111101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001101101011010110100111001111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001101101011010110100111001111001110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111101111011110110011100111001100111001110011101101011010110101101011010110101101100111001110011100111001110011100101100011000111011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111011000110011110110011100111001101101011010110101101011010110101101011010110101101001110011100111100111001110011100111001110010110011101111011111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111011000110011110110011100111001101101011010110101101011010110101101011010110101101001110011100111100111001110011100111001110010110011101111011111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111110111101011000110011001110011100111001100111001110011100111001110110100111001110011100111011010110101101011011001110011100111001110011100101100011001111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001011000110011001110011100111001100111001110011101101011010110101101011010011100111011010110101101011010110101101100111001110011100111001110011100111001100111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111110011100111001011000110011001110011100111001100111001110011101101011010110101101011010011100111011010110101101011010110101101100111001110011100111001110011100111001100111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100100111011010110110011100111001110011100110011101101011011010100111001110110101101011010110101101011010110101101011010110101101100110011100111011010110101101011010110100110110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100100111011010110110011100111001110011100110011101101011011010100111001110110101101011010110101101011010110101101011010110101101100110011100111011010110101101011010110100110110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011011010110100111001110110101101011010011100111001111010110101101010110101101011010011100111001110011100111001110011100111001110011100111011010110101101011010110100111100111001111011111111111111111111111111"),
                ("1111111111111111111111111111111100111001110011001110011101101011010110101101011011010110101101011000110101101010011100111001110011100110100111010110101100001001010011100010011100111011010110101101001110011110011100111001011001111011110111111111111111"),
                ("1111111111111111111111111111111100111001110011001110011101101011010110101101011011010110101101011000110101101010011100111001110011100110100111010110101100001001010011100010011100111011010110101101001110011110011100111001011001111011110111111111111111"),
                ("1111111111111111111111111110011100111001100111001110011101101011010110100111001101001010010100111010110101101011010100111001111010110100100101001010010100111010110101101011010110101001110110101101011010110100111100111001110010110001100111111111111111"),
                ("1111111111111110110001100110011011010110100111100111001100111001110110110101101001001010010100111000100111001110011110101101001001010010100101001010011101010110101101001111000110001101010110101101011010110100111100111001110011111111111111111111111111"),
                ("1111111111111110110001100110011011010110100111100111001100111001110110110101101001001010010100111000100111001110011110101101001001010010100101001010011101010110101101001111000110001101010110101101011010110100111100111001110011111111111111111111111111"),
                ("1111111111111111100111001110011011010110100111100111001110011100110110100111001111010110101101001001110101101011000010010100101001010010100111010110101101010110101101001111000110001101010110101101011010110100111011010110101101111111111111111111111111"),
                ("1111111111111111100111001110011100111001100111001110011100111001111010110101101011010110001100001001010010100101001010000100001001010010100111000110001100011010110100100101001010011101010110101101011010110101101011010110100111100111001111111111111111"),
                ("1111111111111111100111001110011100111001100111001110011100111001111010110101101011010110001100001001010010100101001010000100001001010010100111000110001100011010110100100101001010011101010110101101011010110101101011010110100111100111001111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110100111001101001010010100111010010010100111000010010100101001010000100001001010011100001001010010100101001010011101011000110001001110110101101011010110101101011010110110011100111001111111111111111"),
                ("1111111111111111100111001110011001110011101101001110011100111001111000010010100101001010010100101001110001100001001010000100001000010000100101001010010100111000110001001110110101101011010110101101011010110101101001110011110011100111001111111111111111"),
                ("1111111111111111100111001110011001110011101101001110011100111001111000010010100101001010010100101001110001100001001010000100001000010000100101001010010100111000110001001110110101101011010110101101011010110101101001110011110011100111001111111111111111"),
                ("1111111111111111100111001110011011010110101101011010110100111001111000010010100101001010010100111000010010100101001010000100001000010000100001001010011100001001010011101010110101101001110110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011011010110101101011010110100111001111000010010100101001010010100111000010010100101001010000100001000010000100001001010011100001001010011101010110101101001110110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001101101011010110101101011011010010010100101001010010100101001010000100001000010000100001000010000100001001010011100001001010010100111010110101100011010110101011010110101101100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011001110011100111101011010110101101010011110101101010011110101101001001010000100001000010000100001000010000100001001010011100001001010011100011010110101101001001010011001110011101101100111001011000110001100111111111111111"),
                ("1111111111111111100111001110011001110011100111101011010110101101010011110101101010011110101101001001010000100001000010000100001000010000100001001010011100001001010011100011010110101101001001010011001110011101101100111001011000110001100111111111111111"),
                ("1111111111111111100111001110011011010110110101001110011101101011010110101101011010110110101101001001010010100111000010000100001000010000100001001010011100001001010011001110110101101001111010110101101011010101101100111001111011111111111111111111111111"),
                ("1111111111111111100111001110011001110011110101101011010100111001110011110101101011000010010100101001010010100101001010000100001000010000100001001010011100001001010011101010011100111001110110101101001110011101101001110011110011111111111111111111111111"),
                ("1111111111111111100111001110011001110011110101101011010100111001110011110101101011000010010100101001010010100101001010000100001000010000100001001010011100001001010011101010011100111001110110101101001110011101101001110011110011111111111111111111111111"),
                ("1111111111111111100111001110011001110011110001100011000100111001111010010010100101001010010100111000010010100101000010000100001000010000100101001010010100101001010010100111000110001101010110101101011010110101101001110011110010110001100111111111111111"),
                ("1111111111111111100111001110011001110011100111001110011100111001101001010010100101001010010100111000010010100101001010000100001000010000100101000010000100011000110000100111010110101001110110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011001110011100111001110011100111001101001010010100101001010010100111000010010100101001010000100001000010000100101000010000100011000110000100111010110101001110110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111111111111110011100111001100111011010110100111001101001010010100101001010010100101001010010100101001010000100001000010000100001000010000100001001010011100011010110101001111001110011100111001110011100111001110011111111111111111111111111"),
                ("1111111111111111111111111011001100111001110011001110011101101011010011110101101001001010010100101001010000100001000010000100001000010000100001000010000100111000110001100010011100111001110011100111100111001011000110001100110011111111111111111111111111"),
                ("1111111111111111111111111011001100111001110011001110011101101011010011110101101001001010010100101001010000100001000010000100001000010000100001000010000100111000110001100010011100111001110011100111100111001011000110001100110011111111111111111111111111"),
                ("1111111111111110110001100110011100111001100111011010110101101011010110101101011011010010010100111000010010100101000010000100001000010000100001001010010100101001010011100010011100111101010110101101001110011110010110001100110011100111001111111111111111"),
                ("1111111111111110110001100110011100111001100111011010110101101011010110101101011011010010010100111000010010100101000010000100001000010000100001001010010100101001010011100010011100111101010110101101001110011110010110001100110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010110100111001111010010010100101001010000100001000010000100001000010000100001001010010100101001010011101010110101101001111010110101001110011110011100111001011000110001100111111111111111"),
                ("1111111111111111100111001110011001110011101101011010110101101011010110100111001111000010010100101001010000100001000010000100001000010000100001001010010100101001010011001110110101101001101001010011101011010110010110001100111100110001100111111111111111"),
                ("1111111111111111100111001110011001110011101101011010110101101011010110100111001111000010010100101001010000100001000010000100001000010000100001001010010100101001010011001110110101101001101001010011101011010110010110001100111100110001100111111111111111"),
                ("1111111111111111100111001110011100111001101101011010110101101011010110101101011011010010010100101000010000100001000010000100001000010000100001001010010100101001010011001110110101101011010011100111001110011100110110001100111101110111101111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010110101101011010011010010100101001010010100101000010000100001000010000100001000010000100101001010011101010110101101011011010110100100101001100111100111001011101111011110111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010110101101011010011010010100101001010010100101000010000100001000010000100001000010000100101001010011101010110101101011011010110100100101001100111100111001011101111011110111111111111111"),
                ("1111111111111111100111001110011100111001110011011010110101101011010110101101011010110110101101001001010000100001000010000100001000010000100001000010000100101001010011101010110101101011010011100111101011010100111100111001011000110001100111111111111111"),
                ("1111111111111111111111111110010110001100011001100111001101101011010110101101011010011110101101001001010010100101001010010100101000010000100001000010000100001001010011001110110101101011010011100111011010110110010110001100111111111111111111111111111111"),
                ("1111111111111111111111111110010110001100011001100111001101101011010110101101011010011110101101001001010010100101001010010100101000010000100001000010000100001001010011001110110101101011010011100111011010110110010110001100111111111111111111111111111111"),

                -- 7_explosion_1_1
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111110011100111001110011100111001110010110001100111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011100101100011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111110011100111001110011100111001110010110001100111111111111111110011100111001110011100111001110011100111001110011100111001110011100111001110011100101100011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001110011100111001110011100111001011000110011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0110001100110011100111001110011001110011110011100111001110011100111001100111001110011100111001110110100111001111001101101011010011100111100111001110011011010110101101100111001110011100101100011001111111111111111111111111111111111111111111111111111111"),
                ("0110001100110011100111001110011001110011110011100111001110011100111001100111001110011100111001110110100111001111001101101011010011100111100111001110011011010110101101100111001110011100101100011001111111111111111111111111111111111111111111111111111111"),
                ("0110001100110011001110011101101011010110100111001110011110011100110011100111001111000110101101011010100111001110110101101011010110101101001110011100111001110011100111001111001110011100110011100111100111001111111111111111111111111111111111111111111111"),
                ("1100111001101101011010110101101011010110101101011010110100111001110110100111001111000110101101010011110101101010110101101011010011100111011010011100111100111001110011001110011100111011010110101101100111001111011111111111111111111111111111111111111111"),
                ("1100111001101101011010110101101011010110101101011010110100111001110110100111001111000110101101010011110101101010110101101011010011100111011010011100111100111001110011001110011100111011010110101101100111001111011111111111111111111111111111111111111111"),
                ("1011010110101101011010110101101011010110101101011010110101101011010011100111001110011100111001110110110101101010110100111001110011100111001110011100111100110011100111011010110101101001111001110010110001100011000110001100111101111111111111111111111111"),
                ("1011010110101101011010110101101011010110101101011010110101101011010011100111001110011100111001110110110101101010110100111001110011100111001110011100111100110011100111011010110101101001111001110010110001100011000110001100111101111111111111111111111111"),
                ("1011010110101101011010110101101011010110101101011010110100111001101001010010100111010100111001110110100111001111010110001100011000110000100111010110101011010110101101011010110101101011011001110011100111001110011111011110111101111111111111111111111111"),
                ("1011010110101101011010110101101001110011100111011010110110101101001001010010100101001110101101010110110101101001001010010100101001010010100111010110101001111010110101001110110101101011011001110011100111001110011100111001110011111111111111111111111111"),
                ("1011010110101101011010110101101001110011100111011010110110101101001001010010100101001110101101010110110101101001001010010100101001010010100111010110101001111010110101001110110101101011011001110011100111001110011100111001110011111111111111111111111111"),
                ("1001110011101101001110011110101100011000110101101011010010010100101001010010100101001110001100010110100111001101001010010100101001010011101011010110101101001001010010100111010110101001110011100111100111001110011100111001110011111111111111111111111111"),
                ("1101011010110100100101001010010100101001010010100101001010010100101001010010100101001010010100111010110101101001001010010100101001010010100111000110001101001001010010100111010110101001110110101101001110011100111011010110100111100111001111111111111111"),
                ("1101011010110100100101001010010100101001010010100101001010010100101001010010100101001010010100111010110101101001001010010100101001010010100111000110001101001001010010100111010110101001110110101101001110011100111011010110100111100111001111111111111111"),
                ("0100101001010010100101001010000100101001010011100011000010010100101001110001100011000010010100101001010010100101001110001100001001010011100001001010010100111000110001101011000110001101011010110101001110011100111011010110100111100111001110011111111111"),
                ("0100101001010000100101001010000100001000010000100101001010000100001001010010100101001010010100101001010000100001000010010100111000110000100101001010011101010011100111101011010110101101010011100111011010110100111011010110101101011010110100111111111111"),
                ("0100101001010000100101001010000100001000010000100101001010000100001001010010100101001010010100101001010000100001000010010100111000110000100101001010011101010011100111101011010110101101010011100111011010110100111011010110101101011010110100111111111111"),
                ("0100101001010000100001000010000100001000010000100001000010000100001001010010100101000010010100111000010000100001000010010100101001010010100101001010011100010011100111101010011100111011010110101101011010110101101011010110101101011010110100111111111111"),
                ("0100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100111010110101001110011100111011010110101101011010110100111011010110101101001110011110011111111111"),
                ("0100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100111010110101001110011100111011010110101101011010110100111011010110101101001110011110011111111111"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010011101010011100111001110110101101001110011100111011010110101101100111001011001111111111"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010100101001010011101010011100111001110110101101001110011100111011010110101101100111001011001111111111"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010010100101001010000100001000010000100001000010000100001001010011100001001010010100101001010010100101001010011001110110101101011010110101101001110011110011100111001011001101011010"),
                ("0100001000010000100001000010010100101001010010100101001010000100001000010000100001001010010100101001010010100101001010010100101001010010100111000110001101001001010010100111010110101001110110101101011010110101101001110011110011100111001111101101011010"),
                ("0100001000010000100001000010010100101001010010100101001010000100001000010000100001001010010100101001010010100101001010010100101001010010100111000110001101001001010010100111010110101001110110101101011010110101101001110011110011100111001111101101011010"),
                ("0100001000010010100101001010010100101001010010100101001010010100101000010000100001001110001100011000110001100011000110001100001001010010100111000110001101011010110100100111000110001001110110101101011010110101101100111001110011100111001110011001110011"),
                ("0100101001010010100101001010010100101001010010100101001110001100001001110001100001001010010100101001010010100101001010010100111000110000100111010110101011010110101101101001001010011001110110101101011010110110011100111001110011100111001111111101011010"),
                ("0100101001010010100101001010010100101001010010100101001110001100001001110001100001001010010100101001010010100101001010010100111000110000100111010110101011010110101101101001001010011001110110101101011010110110011100111001110011100111001111111101011010"),
                ("1001110011110101101011010100111001110011110101100011000110001100011000010010100101001110101101010011110001100001001110101101010011100111101001001010011001110011100111101011000110001001111001110011100111001110011100111001110011111111111111111001110011"),
                ("1011010110101101011010110101101011010110101101001110011100111001111010110101101011000100111001110110110101101011010101101011010110101101100001001010011100011000110001101010011100111001110011100111100111001110011100111001011001111111111111111001110011"),
                ("1011010110101101011010110101101011010110101101001110011100111001111010110101101011000100111001110110110101101011010101101011010110101101100001001010011100011000110001101010011100111001110011100111100111001110011100111001011001111111111111111001110011"),
                ("1011010110101101011010110101101001110011100111101011010100111001110011100111001111010100111001110011110101101011000100111001110110101101001111010110101101011010110101001110110101101011010110101101100111001110010110001100011101111111111111111001110011"),
                ("1001110011100111101011010100110100101001110101011010110100111001111001101101011010110101101011011010010010100111010101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001011001110111101111111111111111111111100111001"),
                ("1001110011100111101011010100110100101001110101011010110100111001111001101101011010110101101011011010010010100111010101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001011001110111101111111111111111111111100111001"),
                ("1011010110110100100101001100111101011010100111001110011110011100111001101101011010110100111001111010100111001110110101101011010110101101011010110101101011010110101101011010011100111011010110101101100111001111101111111111111111111111111111111111111111"),
                ("1011010110110100100101001100111101011010100111001110011110011100111001101101011010110100111001111010100111001110110101101011010110101101011010110101101011010110101101011010011100111011010110101101100111001111101111111111111111111111111111111111111111"),
                ("1100111001100111001110011100111100111001110011100111001011000110011001100111001110110101101011010110101101011010110100111001110110101101011010110101101001110011100111001111001110011001110011100111001110011111111111111111111111111111111111111111111111"),
                ("0110001100110011100111001011000110001100110010110001100011000110011001110011100110011100111001111001110011100111001110011100110011100111011010110101101011011001110011100111001110011100101100011001111111111111111111111111111111111111111111111111111111"),
                ("0110001100110011100111001011000110001100110010110001100011000110011001110011100110011100111001111001110011100111001110011100110011100111011010110101101011011001110011100111001110011100101100011001111111111111111111111111111111111111111111111111111111"),
                ("1111111111011000111001110111101111011110011001100111001110011100111001110011100111001110011100111101011000110011001110011100111001110011100110011100111011011001110011100101100011001110111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111011001111011110111010110001100011001100111001111111111111111110011100101100111111111111111011000110011001110011100111001110011100111001110011111111111111110110011110111101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111011001111011110111010110001100011001100111001111111111111111110011100101100111111111111111011000110011001110011100111001110011100111001110011111111111111110110011110111101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_1_2
                ("1111111111111111111111111111110110001100110011011010110100111001110110101101011010011010010100101000010000100001000010000100001001010010100101001010010100111010110101001110110101101011010110101101100111001011000110001100110011111111111111111111111111"),
                ("1111111111111111111111111111110110001100110011011010110100111001110110101101011010011010010100101000010000100001000010000100001001010010100101001010010100111010110101001110110101101011010110101101100111001011000110001100110011111111111111111111111111"),
                ("1111111111111110110001100011001100111001100111101011010100111001110110101101011011010010010100101001010000100001000010000100001000010000100001000010000100111010110101011010110101101011010110101101011010110110011100111001110011100111001111111111111111"),
                ("1111111111111111111011110011101100111001100110100101001110101101010110101101011011010010010100101001010000100001000010000100001000010000100001001010010100101001010011001110110101101011010110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111111011110011101100111001100110100101001110101101010110101101011011010010010100101001010000100001000010000100001000010000100001001010010100101001010011001110110101101011010110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111110111101111100110001100100111001110011100111001110110101101011010011010010100101001010010100101000010000100001000010000100001000010000100001001010011101010110101101011010110101101011010110101101100111001110011100111001111111111111111"),
                ("1111111111111110110001100111100110001100110011101011010010010100110011101101011010011010010100101001010010100101000010000100001000010000100001000010000100101001010011100010011100111011010110101101011010110101101001110011110011100111001111111111111111"),
                ("1111111111111110110001100111100110001100110011101011010010010100110011101101011010011010010100101001010010100101000010000100001000010000100001000010000100101001010011100010011100111011010110101101011010110101101001110011110011100111001111111111111111"),
                ("1111111111111110110001100011001100111001110011001110011110101101010011101101011011010010010100101001010010100101000010000100001000010000100001000010000100101001010011101010011100111011010110101101011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001110010110001100110011001110011101101011011010100111001111000010010100101001010010100101000010000100001000010000100001001010011100001001010011101010110101101011010110101101011010110100111100111001110010110001100111111111111111"),
                ("1111111111111111100111001110010110001100110011001110011101101011011010100111001111000010010100101001010010100101000010000100001000010000100001001010011100001001010011101010110101101011010110101101011010110100111100111001110010110001100111111111111111"),
                ("1111111111111111111111111110010110001100011001100111001100111001110011100111001111000110001100001001010000100001000010000100001000010000100001000010000100101001010010100111010110101001110110101101001110011110011100111001011001111111111111111111111111"),
                ("1111111111111111111111111110010110001100011001100111001100111001110011100111001111000110001100001001010000100001000010000100001000010000100001000010000100101001010010100111010110101001110110101101001110011110011100111001011001111111111111111111111111"),
                ("1111111111111111111111111110011100111001110011100111001110011100110011110101101011000010010100101000010000100001000010000100001000010000100101001010010100101001010010100101001010010100110011100111011010110100111100111001110011111111111111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010011110101101001001110001100001000010000100001001010000100001000010000100101001010011100001001010010100101001010010100110011100111001110011100111001110011110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010011110101101001001110001100001000010000100001001010000100001000010000100101001010011100001001010010100101001010010100110011100111001110011100111001110011110011100111001111111111111111"),
                ("1111111111111110110001100110011001110011101101011010110101101011011010110001100001001010010100101001010010100101001010000100001000010000100001001010011100001001010010100101001010011101010011100111100011000110001001110011110011100111001111111111111111"),
                ("1111111111111111111111111110011001110011101101001110011101101011010011100111001111010010010100111000010010100101000010000100001000010000100101001010010100101001010011100011010110101001110011100111101011010110101001110011110011100111001111111111111111"),
                ("1111111111111111111111111110011001110011101101001110011101101011010011100111001111010010010100111000010010100101000010000100001000010000100101001010010100101001010011100011010110101001110011100111101011010110101001110011110011100111001111111111111111"),
                ("1111111111111111111111111111011100111001101101101011010110101101010011101101011010011010010100111000010010100101000010000100001000010001100001001010010100111010110101011010110101101011010110101101001110011110101011010110110011100111001111111111111111"),
                ("1111111111111110110001100011001100111001101101001110011010010100111010110101101011000010010100111000010010100101000010000100001000010000100001000010000100111010110101001111010110101001111010110101101011010100111001110011110011100111001111111111111111"),
                ("1111111111111110110001100011001100111001101101001110011010010100111010110101101011000010010100111000010010100101000010000100001000010000100001000010000100111010110101001111010110101001111010110101101011010100111001110011110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001101101011010110110101101011000110101101001001010010100111000010010100101000010000100001000010000100001000010000100101001010010100101001010011101010110101101011010110101101100111001110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010011101101011011010010010100111000010010100101000010000100001000010000100101001010011100001001010010100101001010011100010011100111011010110101101011010110110011100111001111111111111111"),
                ("1111111111111111100111001110011100111001100111011010110101101011010011101101011011010010010100111000010010100101000010000100001000010000100101001010011100001001010010100101001010011100010011100111011010110101101011010110110011100111001111111111111111"),
                ("1111111111111111100111001110011001110011101101011010110101101011010110101101011010011110001100001001010010100101001010000100001000010000100111000110000100101001010010100101001010011100010011100111001110011101101001110011110011100111001111111111111111"),
                ("1111111111111111100111001110011001110011101101011010110101101011010110101101011010011110001100001001010010100101001010000100001000010000100111000110000100101001010010100101001010011100010011100111001110011101101001110011110011100111001111111111111111"),
                ("1111111111111111100111001110011011010110101101011010110101101011010011110001100011010010010100101001010010100111000010010100101000010000100101001010011100001001010011101001001010010100110011100111011010110100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001100111011010110101101011010110101101011011010010010100101001110101101011000110001100001001010010100101000010000100101001010010100111000110001101011010110101101010011100111001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111100111001100111011010110101101011010110101101011011010010010100101001110101101011000110001100001001010010100101000010000100101001010010100111000110001101011010110101101010011100111001110011100111100111001110011100111001111111111111111"),
                ("1111111111111111111111111101101011010110100111011010110101101011011010110001100010011101101011011010110101101001001010010100101001010011100011010110100100111010110101101010011100111011011001110011100111001100111011010110110011100111001111111111111111"),
                ("1111111111111111111111111110011100111001100111011010110101101011011010110001100010011101101011011010010010100101001010010100111010110101001110011100111100001001010010100111010110101011010011100111100111001100111011010110110010110001100111111111111111"),
                ("1111111111111111111111111110011100111001100111011010110101101011011010110001100010011101101011011010010010100101001010010100111010110101001110011100111100001001010010100111010110101011010011100111100111001100111011010110110010110001100111111111111111"),
                ("1111111111111110110001100110011100111001100111011010110101101011010011110101101011010110101101001001010010100101001110101101010011100111101011010110101101001001010010100110011100111011010110101101001110011100111100111001110011111111111111111111111111"),
                ("1111111111111111111011110011001100111001110011001110011101101011010110100111001111000010010100111000110101101001001100111001110011100111001111010110101100011010110101101010110101101011010110101101001110011110011100111001111111111111111111111111111111"),
                ("1111111111111111111011110011001100111001110011001110011101101011010110100111001111000010010100111000110101101001001100111001110011100111001111010110101100011010110101101010110101101011010110101101001110011110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111011100111001100111011010110101101011010110100111001110011100111001110011100111001110011100111001110110101101011011010110101101010011100111001110110101101011010011100111011010110110011100111001111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100100111011010110101101011010110100111001111001101101011010110101101011010110101101011010110101101011010011100111101010110101101001111001110011100111001110011011010110100110110001100111111111111111111111111111111"),
                ("1111111111111111111111111111110110001100100111011010110101101011010110100111001111001101101011010110101101011010110101101011010110101101011010011100111101010110101101001111001110011100111001110011011010110100110110001100111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111100111100111001110011100111001110011100111001101101011010110101101011010110100111001110110101101011010110101101001110011100111100111001110011100101100011001100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111100111100111001110011100111001110011100111001101101011010110101101011010110100111001110110101101011010110101101001110011100111100111001110011100101100011001100111001110011111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110011000110011001110011100111001110011100110110101101011010110100111001110011100111011010011100111001110011100111100111001110011100101100011001110111101111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111011110101100110011100111001110011100111001100111001110011101101011010110101101011010110101101011010110101101100111001110011111001100011001111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111011110101100110011100111001110011100111001100111001110011101101011010110101101011010110101101011010110101101100111001110011111001100011001111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111101110011000110011001110011100111001110011100111001101101011010110101101011010110101101001110011100111100111001110011111011110111101111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011100110011100111011010110101101100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011100110011100111011010110101101100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101111001100011000110011001110011001110011100111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111110011100110011100111001110011110101101010011110101101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111110011100110011100111001110011110101101010011110101101011010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_1_3
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111101111001100111111111111111110011100111001110011100111001110011100101100011001111111111111110110011001110011111111111111111100111001011000110001100111011111011110011001111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111101111001100111111111111111110011100111001110011100111001110011100101100011001111111111111110110011001110011111111111111111100111001011000110001100111011111011110011001111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111101011000110011001110011100110110100111001111001110011100111001110011100101100011001110111001110011100111001110011100111001110011100111001011001111011110111100111001110011001111111111"),
                ("1111111111111111111111111111111111111111111111111111111011000110011001110011100111001110011100110110101101011010110100111001111001110011100111001110011100110011100111001111001110011100101100011000110001100110010110001100011001100111001110010110001100"),
                ("1111111111111111111111111111111111111111111111111111111011000110011001110011100111001110011100110110101101011010110100111001111001110011100111001110011100110011100111001111001110011100101100011000110001100110010110001100011001100111001110010110001100"),
                ("1111111111111111111111111111111111111111111111001110011100111001110011110011100110011100111001110011101101011010110101101011010011100111011010110101101011010110101101011010011100111100101100011001100111001110011100111001100111001110011100111100111001"),
                ("1111111111111111111111111111111111111111111101100111001101101011010110100111001110110101101011010110101101011010110101101011010110101101011010011100111101010011100111011010110101101100111001110011001110011100111101011010100110100101001110101011010110"),
                ("1111111111111111111111111111111111111111111101100111001101101011010110100111001110110101101011010110101101011010110101101011010110101101011010011100111101010011100111011010110101101100111001110011001110011100111101011010100110100101001110101011010110"),
                ("1100111001111111111111111111111110111101011001100111001101101011010110101101011010110101101011010110101101011010110101101011010110101101101001001010011101010110101101011010110101101100110011100111011010110110100100101001100111101011010100111001110011"),
                ("1100111001111111111111111111111110111101011001100111001101101011010110101101011010110101101011010110101101011010110101101011010110101101101001001010011101010110101101011010110101101100110011100111011010110110100100101001100111101011010100111001110011"),
                ("1001110011111111111111111011100110001100110011100111001101101011010110101101011010011110101101011010110101101010011101101011010011100111100011010110101001110011100111101010011100111001110011100111101011010100111001110011101101011010110101101011010110"),
                ("1001110011111111111111111011001100111001110011100111001100111001110011100111001111010110001100011000010010100111000101101011010110101101101011010110101011010011100111100011010110101101010011100111001110011101101011010110101101011010110101101011010110"),
                ("1001110011111111111111111011001100111001110011100111001100111001110011100111001111010110001100011000010010100111000101101011010110101101101011010110101011010011100111100011010110101101010011100111001110011101101011010110101101011010110101101011010110"),
                ("1001110011111111111111111110011100111001110011100111001110011100110011110001100011010100111001110011010010100111010100111001111010110100100111000110001001111010110100100101001010011100011000110001100011000110101001110011100111101011010110101001110011"),
                ("1101011010111111100111001110011100111001110011011010110101101011010011010010100111010101101011010110110101101001001110001100001001010010100101001010010100101001010010100111000110000100111000110000100101001010010100101001010010100101001010010100101001"),
                ("1101011010111111100111001110011100111001110011011010110101101011010011010010100111010101101011010110110101101001001110001100001001010010100101001010010100101001010010100111000110000100111000110000100101001010010100101001010010100101001010010100101001"),
                ("1001110011110011100111001110011100111001101101011010110101101011010011110001100001001110101101011010110001100001001010010100111000110001100011000110001100011000110000100101000010000100001001010010100101001010010100101001010010100101001010010100001000"),
                ("1101011010111101100111001110011001110011101101011010110101101011010011110101101001001010010100111010110001100001001010010100101001010010100101001010010100101001010010100101000010000100001000010000100101001010010100101001010010100001000010000100001000"),
                ("1101011010111101100111001110011001110011101101011010110101101011010011110101101001001010010100111010110001100001001010010100101001010010100101001010010100101001010010100101000010000100001000010000100101001010010100101001010010100001000010000100001000"),
                ("1101011010011001100111001110011001110011101101011010110101101011010011010010100101001010010100101001010010100111000010010100101000010000100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001000010000100001000"),
                ("1111111111011001100111001101101011010110100111001110011101101011010011100111001111010010010100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("1111111111011001100111001101101011010110100111001110011101101011010011100111001111010010010100101001010010100101001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("1111111111110011001110011101101011010110100111011010110101101011010110100111001110011110101101001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001"),
                ("1111111111110011001110011101101011010110100111011010110101101011010110100111001110011110101101001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001"),
                ("1111111111100111011010110101101011010110101101011010110101101011010110100111001111010100111001111000010010100101001010010100101001010010100001000010001100001001010010100001001010010100101000010000100001000010000100001000010000100001000010000100101001"),
                ("1111111111100111011010110101101011010110100111011010110100111001111010110101101011010100111001111010010010100101001110001100001001010010100001000010000100101001010010100101001010010100101000010000100101001010000100001000010000100101001010000100101001"),
                ("1111111111100111011010110101101011010110100111011010110100111001111010110101101011010100111001111010010010100101001110001100001001010010100001000010000100101001010010100101001010010100101000010000100101001010000100001000010000100101001010000100101001"),
                ("1111111111110011100111001100111011010110100111001110011110101101011010110001100011010110001100001001010010100111000010010100111000110000100101001010010100101001010011100011000110000100101001010011100011000010010100101001010000100101001010010100101001"),
                ("1111111111111111100111001100111011010110100111001110011101101011010011110101101001001010010100111010110001100001001010010100101001010010100111010110101101001001010010100101001010010100101001010010100101001010010100101001010010100101001110101101011010"),
                ("1111111111111111100111001100111011010110100111001110011101101011010011110101101001001010010100111010110001100001001010010100101001010010100111010110101101001001010010100101001010010100101001010010100101001010010100101001010010100101001110101101011010"),
                ("1111111111111111111111111110011100111001110011100111001100111001110011110101101001001010010100111010110101101011010010010100101001010010100110011100111011011000110000100101001010010100101001010011101011010110101100011000110101001110011101101001110011"),
                ("1111111111111111111111111110011100111001110011100111001110011100110110101101011010011110101101010011110101101001001010010100101001010010100111010110101011011010110100100101001010010100111010110101011010110100111001110011101101011010110101101011010110"),
                ("1111111111111111111111111110011100111001110011100111001110011100110110101101011010011110101101010011110101101001001010010100101001010010100111010110101011011010110100100101001010010100111010110101011010110100111001110011101101011010110101101011010110"),
                ("1111111111111111111111111111101111011110110011100111001110011100110110101101011010110101101011010110110101101001001110001100011000110001101010011100111011010011100111101001001010010100110011100111011010110101101011010110101101011010110101101011010110"),
                ("1111111111111111111111111111100110001100011000110001100110011100110011101101011010110100111001111001100111001110011100111001110011100111011011010110101011010011100111001110011100111001110110101101011010110101101011010110101101011010110101101011010110"),
                ("1111111111111111111111111111100110001100011000110001100110011100110011101101011010110100111001111001100111001110011100111001110011100111011011010110101011010011100111001110011100111001110110101101011010110101101011010110101101011010110101101011010110"),
                ("1111111111111111111111111111111111111111111011100111001101101011010110100111001110011110011100111001100111001110110100111001110110101101011011010110101001111010110101100010011100111011010011100111011010110101101011010110101101011010110101101100111001"),
                ("1111111111111111111111111111111111111111111011100111001101101011010110100111001110011110011100111001100111001110110100111001110110101101011011010110101001111010110101100010011100111011010011100111011010110101101011010110101101011010110101101100111001"),
                ("1111111111111111111111111111111111111111111111100111001100111001111001110011100110011100111001110011100111001110011101101011010110101101011010011100111101011010110101100010011100111001111001110011001110011100111011010110101101001110011110010110001100"),
                ("1111111111111111111111111111111111111111111111111111111011000110011001110011100111001101101011010110110011100111001100111001110110101101100110011100111011010011100111001110011100111100111001110011100111001110011001110011110011100111001110010110001100"),
                ("1111111111111111111111111111111111111111111111111111111011000110011001110011100111001101101011010110110011100111001100111001110110101101100110011100111011010011100111001110011100111100111001110011100111001110011001110011110011100111001110010110001100"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100101100011001100111001110011100111001110011100111001110011100111001"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000110011001110011100111001110011100111001110011100111001110011100111001110011100111001110011111111111111110110001100110011100111001110011100111001110011111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000110011001110011100111001110011100111001110011100111001110011100111001110011100111001110011111111111111110110001100110011100111001110011100111001110011111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_2_0
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001111101111001100011000110011000110000110011110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001111101111001100011000110011000110000110011110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100110011100111001110011100110011100111011010110101101100101100011000110011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111011100111001100011000110001100110011100111001110011100110011100111011010110101101001111001110011100111001110011111011110111101111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111011100111001100011000110001100110011100111001110011100110011100111011010110101101001111001110011100111001110011111011110111101111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111110011000110011001100111001111001110011100111001110011100110011100111011010110101101011010110101101001111001110010110001100011001100111001111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111101111011110110011100110011101101011010110101101011010110101101011010110101101011010011100111001110110101101001111001110011100111001110011100111001111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111101111011110110011100110011101101011010110101101011010110101101011010110101101011010011100111001110110101101001111001110011100111001110011100111001111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111110111001110111101111011001110011100110110101101011010110100111001110011100111001110110101101011010011100111100010011100111011010110101101100111001110011100111001011000110001100111111111111111111111111111111"),
                ("1111111111111111111111111100111100111001011000111001110110011100111001110011100110110101101011010110100111001110110100111001110011100111001111000110000100001000010001100010011100111011010110101101011010110101100110001100011001111111111111111111111111"),
                ("1111111111111111111111111100111100111001011000111001110110011100111001110011100110110101101011010110100111001110110100111001110011100111001111000110000100001000010001100010011100111011010110101101011010110101100110001100011001111111111111111111111111"),
                ("1111111111111111111111111111100110001100110010110001100110011100110011110011100110110101101011011010100111001110110110101101011000110001100001001010010100001000010001100010110101101011010110101101011010110101101001110011011001111011110111111111111111"),
                ("1111111111111111111111111111100110001100110010110001100110011100110011110011100110110101101011011010100111001110110110101101011000110001100001001010010100001000010001100010110101101011010110101101011010110101101001110011011001111011110111111111111111"),
                ("1111111111111111111111111111111110111101011001111011110011000110010110100111001110011110101101001001110001100011010110001100001001010010100101001010010100001000010000100111010110101011010110101101011010110100111100111001111010111001110111101111111111"),
                ("1111111111111111111111111111111100111001110010110001100110011100110110101101011010110100111001101001010010100101001010010100111000110000100101001010010100001000010000100011000110001001110110101101011010110100111100111001011000110001100111101111111111"),
                ("1111111111111111111111111111111100111001110010110001100110011100110110101101011010110100111001101001010010100101001010010100111000110000100101001010010100001000010000100011000110001001110110101101011010110100111100111001011000110001100111101111111111"),
                ("1111111111111111111111111011001100111001101101001110011100111001110110101101011010110010010100101001010000100001000010000100001001010010100101000010000100001000010000100011010110101001110110101101011010110101101100111001110010110001100111101111111111"),
                ("1111111111111111111111111110011100111001101101011010110101101011010110101101011010011010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100111010110101011010110101101001110011110011100111001011001111111111"),
                ("1111111111111111111111111110011100111001101101011010110101101011010110101101011010011010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100111010110101011010110101101001110011110011100111001011001111111111"),
                ("1111111111111111111111111110011001110011100111011010110101101011010110101101011010011010010100101000010010100101000010000100001000010000100001000010000100001000010000100011000110000100111010110101011010110101101011010110100111001110011110011111111111"),
                ("1111111111111111111111111110011001110011110011001110011100111001110011101101011010011010010100101000010000100001001010000100001000010000100001000010000100001001010010100101001010010100111010110101001110011100111100111001100111100111001110011111111111"),
                ("1111111111111111111111111110011001110011110011001110011100111001110011101101011010011010010100101000010000100001001010000100001000010000100001000010000100001001010010100101001010010100111010110101001110011100111100111001100111100111001110011111111111"),
                ("1111111111111111111111111110011100111001110011100111001100111001110011100111001111010010010100101000010010100101000010010100101000010000100001000010000100101001010010100001000010000100111010110101101011010110101101011010110011100111001110011111111111"),
                ("1111111111111111100111001110011100111001110011100111001101101011010110110101101001001110001100011000010010100101000010000100001000010001011101000010000100001001010010100001000010000100110011100111101011010110101001110011100111100111001110011111111111"),
                ("1111111111111111100111001110011100111001110011100111001101101011010110110101101001001110001100011000010010100101000010000100001000010001011101000010000100001001010010100001000010000100110011100111101011010110101001110011100111100111001110011111111111"),
                ("1111111111011001100111001110011100111001110011001110011100111001111010110001100001001010010100101001010000100001000010000100010111101110000110111101110100001000010000100001000010001001110110101101001110011100111011010110110010110001100111101111111111"),
                ("1111111111011001100111001110011100111001110011001110011100111001111010110001100001001010010100101001010000100001000010000100010111101110000110111101110100001000010000100001000010001001110110101101001110011100111011010110110010110001100111101111111111"),
                ("1111111111110011100111001100111100111001100111001110011110101101001001010010100101000010000100011000010000100001000010000100001000010001011100001000011011101000010000100101001010011101010011100111001110011100111001110011011000111001110111101111111111"),
                ("1111111111110011100111001101101011010110101101011010110110101101001001010010100101000010010100101001010000100001000110111101110111101111011100001000011011101000010000100001001010011101010011100111001110011100111011010110110010111001110111101111111111"),
                ("1111111111110011100111001101101011010110101101011010110110101101001001010010100101000010010100101001010000100001000110111101110111101111011100001000011011101000010000100001001010011101010011100111001110011100111011010110110010111001110111101111111111"),
                ("1111111111111011110111101110011001110011100111001110011100111001110011110101101001001010000100001000010000100001000000010000110111101110100011011110111101101000010000100101001010011100001001010010100101001100111001110011110010110001100111101111111111"),
                ("1111111111111111111011110011001001110011010010100101001110101101010011110101101001000010000100001000010000100001000000010000110111101110100001000010000100001001010011100001001010010100001000010000100101001100111011010110110010110001100011101111111111"),
                ("1111111111111111111011110011001001110011010010100101001110101101010011110101101001000010000100001000010000100001000000010000110111101110100001000010000100001001010011100001001010010100001000010000100101001100111011010110110010110001100011101111111111"),
                ("1111111111111111111111111011001100111001110101101011010110101101011010110101101001001010000100001000010000100001000101111011111011110110100001000010000100001000010000100001000010000100001000010000100101001100111001110011110011110111101111101111111111"),
                ("1111111111111111111111111011001100111001101101011010110101101011010110110001100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010011101011010100111100111001111010111001110111111111111111"),
                ("1111111111111111111111111011001100111001101101011010110101101011010110110001100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010011101011010100111100111001111010111001110111111111111111"),
                ("1111111111111111111011110011001100111001101101001110011110101101010011010010100101000010000100001000010000100001000010000100001000010001101111011110110100001000010000100101001010010100011000110000100101001100110110001100011101111011110111111111111111"),
                ("1111111111111101110111101110011011010110101101001110011110101101001001010000100001000010000100001000010000100001000010000100011011110110000100001000011011101000010000100111010110101100011010110101101011010100111100111001110011111011110111101111111111"),
                ("1111111111111101110111101110011011010110101101001110011110101101001001010000100001000010000100001000010000100001000010000100011011110110000100001000011011101000010000100111010110101100011010110101101011010100111100111001110011111011110111101111111111"),
                ("1111111111111100110001100110011001110011101101011010110100111001111000010010100101000010000100001000010000100010111110111101110111101110000100001000010000101000010000100111000110000100111010110101101011010100111011010110110011111011110111101111111111"),
                ("1111111111111100110001100110011001110011101101011010110100111001111000010010100101000010000100001000010000100010111110111101110111101110000100001000010000101000010000100111000110000100111010110101101011010100111011010110110011111011110111101111111111"),
                ("1111111111111101111011110011001100111001101101011010110100111001101001010010100101001010000100001000010000100011011101111011100001000011011110111101110000110111101110100010011100111001110011100110100101001100111011010110100111100111001111101111111111"),
                ("1111111111110011100111001110011011010110101101011010110100111001101001010010100101001010000100001000010000100010111101111011110111101110100010111101110000111011110110100011000110001101010011100111001110011101101100111001110011100111001011001111111111"),
                ("1111111111110011100111001110011011010110101101011010110100111001101001010010100101001010000100001000010000100010111101111011110111101110100010111101110000111011110110100011000110001101010011100111001110011101101100111001110011100111001011001111111111"),
                ("1111111111111111100111001110011100111001100111101011010100111001111010010010100101001010000100001000010000100011011101111011100001000010000100001000011011101000010000100111000110000100111000110001011010110101101001110011110011100111001110011111111111"),
                ("1111111111111111110111101011001111011110110011001110011101101011011010010010100111000010000100001000010000100011011101111011110111101111011110111101110000110111101110100010011100111001110011100111011010110101101001110011110011100111001110011111111111"),
                ("1111111111111111110111101011001111011110110011001110011101101011011010010010100111000010000100001000010000100011011101111011110111101111011110111101110000110111101110100010011100111001110011100111011010110101101001110011110011100111001110011111111111"),
                ("1111111111011101111011110110011100111001100111101011010100111001111010010010100101001110001100001001010000100010111101111011100001000010000100001000011011111011110110100001001010011101011010110101011010110101101001110011110011100111001011001111111111"),
                ("1111111111011001100111001011001111011110110011001110011101101011011010010010100111000110001100001001010000100011011110111101110111101110000110111101111101101000010000100001000010000100110011100111011010110101101001110011110011100111001011101111111111"),
                ("1111111111011001100111001011001111011110110011001110011101101011011010010010100111000110001100001001010000100011011110111101110111101110000110111101111101101000010000100001000010000100110011100111011010110101101001110011110011100111001011101111111111"),

                -- 7_explosion_2_1
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0110001100011101111111111111111100111001111101111011110111101111011111111111111111111111111111111101110011100111001011000110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001111101110111101110011100111001111100110001100111011110111110111111111111111111101111011101110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001111101110111101110011100111001111100110001100111011110111110111111111111111111101111011101110011100111001110011100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("0110001100110010110001100110011100111001011001100111001110011100101100011000110001100011000110011001101101011010011110011100111001110011100111001110011100111001110010110011111111111111111110111101001110011111111111111111111111111111111111111111111111"),
                ("1111011110110011111011110110011011010110110011001110011101101011011001110011100111001100111001110011101101011011001110011100111001110011100110011100111001111001110011100111001110011110101100011001100111001111111111111111111111111111111111111111111111"),
                ("1111011110110011111011110110011011010110110011001110011101101011011001110011100111001100111001110011101101011011001110011100111001110011100110011100111001111001110011100111001110011110101100011001100111001111111111111111111111111111111111111111111111"),
                ("1100111001100111100111001100111011010110101101011010110101101011010110101101011011010010010100110011101101011010011110011100111001110011100111001110011001110110101101011011001110010110011001110010110001100111111111111111111111111111111111111111111111"),
                ("1001110011110101001110011110101011010110101101011010110100111001110011101101011011010010010100110011101101011010011100111001111001110011100110011100111011010110101101001101100011001111001100011000111001110011101111111111111111111111111111111111111111"),
                ("1001110011110101001110011110101011010110101101011010110100111001110011101101011011010010010100110011101101011010011100111001111001110011100110011100111011010110101101001101100011001111001100011000111001110011101111111111111111111111111111111111111111"),
                ("1011010110100111011010110100111001110011100111001110011110101101011010101101011011010110101101010011110101101011010100111001110110101101001110011100111011010110101101001111001110010110011001110011100111001111101111011110111111111111111111111111111111"),
                ("1011010110100111011010110100111001110011100111001110011110101101011010101101011011010110101101010011110101101011010100111001110110101101001110011100111011010110101101001111001110010110011001110011100111001111101111011110111111111111111111111111111111"),
                ("1101011010110101101011010110100100101001010011100011000010010100110011101101011011010100111001110011010010100101001110101101010110101101001110011100111011010110101101011010110101101011010011100111100111001110011111011110111101111111111111111111111111"),
                ("0100101001010010100101001010010100101001010010100101001010000100001001110001100011010110101101011010010010100101001110001100011010110101001110110101101011010110101101011010110101101001111001110011100111001110011100111001011000111001110111111111111111"),
                ("0100101001010010100101001010010100101001010010100101001010000100001001110001100011010110101101011010010010100101001110001100011010110101001110110101101011010110101101011010110101101001111001110011100111001110011100111001011000111001110111111111111111"),
                ("1100011000010011100011000010010100101001010010100001000010000100001000010000100001001010000100001001010000100001000010010100101001010011101010011100111001110011100111011010110101101001110110101101011010110101101001110011110010110001100111111111111111"),
                ("1100011000110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010100101000010010100111000110000100101001010010100101000010000100110011100111101010110101101011010110101101011010110100110110001100111111111111111"),
                ("1100011000110000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010100101000010010100111000110000100101001010010100101000010000100110011100111101010110101101011010110101101011010110100110110001100111111111111111"),
                ("0100101001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010100111000010010100111000110000100001000010000100001000010000100101001010010100111010110101011010110101101011010110110010110001100011001111111111"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100101000010000100001001010011100010011100111001110011100111011010110110011100111001110011100111001"),
                ("0100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100101000010000100001001010011100010011100111001110011100111011010110110011100111001110011100111001"),
                ("1101111011101111101111011110111011110111110111011110111010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100001000010000100001001010011101010110101101011010110100111011010110110011100111001110011100111001"),
                ("1101111011101111011110111101111011110111101111101111011010000100001000010000100010111000010000100001110111101101000010000100001000010000100101000010000100001000010000100001001010011100011010110101001110011100111011010110110011100111001110011111011110"),
                ("1101111011101111011110111101111011110111101111101111011010000100001000010000100010111000010000100001110111101101000010000100001000010000100101000010000100001000010000100001001010011100011010110101001110011100111011010110110011100111001110011111011110"),
                ("1011110111000011011110111000011011110111000011011110111110111101101000010000100011011101111011110111101111011101000101111011101000010000100001000010000100001000010000100111000110000100111000110001001110011101101011010110100111001110011100110110001100"),
                ("1011110111000011011110111000011011110111000011011110111110111101101000010000100011011101111011110111101111011101000101111011101000010000100001000010000100001000010000100111000110000100111000110001001110011101101011010110100111001110011100110110001100"),
                ("0000100001000011011110111000010100001000101110000100001000010000111011010000100001000010000100001000101111011110111000010000110111101110100001000010000100001000010000100101001010010100111000110001001110011101101011010110101101011010110101100110001100"),
                ("1011110111000011011110111000011011110111101110000100001000010000111011010000100001000010000100011011000010000100001101111011101000010000100001000010000100001000010000100001001010010100101001010011100011000100111001110011101101011010110101101100011000"),
                ("1011110111000011011110111000011011110111101110000100001000010000111011010000100001000010000100011011000010000100001101111011101000010000100001000010000100001000010000100001001010010100101001010011100011000100111001110011101101011010110101101100011000"),
                ("1101111011101110000100001101110000100001000010000100001101111011101000010000100001000010000100011011101111011110111010000100001000010000100101000010000100001000010000100001000010000100001000010000100001000110001001110011101101001110011110010110001100"),
                ("0100001000110111011110111010001101111011101110100001000010000100001000010000100001000010010100101000010000100001000010000100001001010010100101001010010100001000010000100001000010000100001000010000100001000100111011010110101101100111001011001111011110"),
                ("0100001000110111011110111010001101111011101110100001000010000100001000010000100001000010010100101000010000100001000010000100001001010010100101001010010100001000010000100001000010000100001000010000100001000100111011010110101101100111001011001111011110"),
                ("0100001000010000100001000010010100001000010000100101001010010100101001010000100001000110001100001001010000100001001010000100001000010000100001001010010100001000010000100001000010000100111000110001100011000101101001110011100111100111001011001111111111"),
                ("0100001000010011001110011110001100011000100111100011000110101101001001010000100001000010010100101001010010100101001010000100001000010000100001001010011100001001010011101011000110001101010110101101001110011101101100111001110011100111001111111111111111"),
                ("0100001000010011001110011110001100011000100111100011000110101101001001010000100001000010010100101001010010100101001010000100001000010000100001001010011100001001010011101011000110001101010110101101001110011101101100111001110011100111001111111111111111"),
                ("0100101001110101001110011010011101011010100110100101001110001100001000010000100001000010000100011000110101101011010100111001101001010010100101001010010100101001010011001110011100111011010110101101011010110110011100111001011001111011110111111111111111"),
                ("1001110011110101001110011110001001110011100111101011010110101101011000010010100101000010000100001001100111001110011101101011010011100111101011010110101101011010110101011010110101101011010110101101011010110110011100111001011001111011110111111111111111"),
                ("1001110011110101001110011110001001110011100111101011010110101101011000010010100101000010000100001001100111001110011101101011010011100111101011010110101101011010110101011010110101101011010110101101011010110110011100111001011001111011110111111111111111"),
                ("1011010110101101011010110101101001110011010011101011010110101101001001110101101001001010010100101001100111001110011100111001111010110101101010011100111011010110101101011010110101101011010110101101011010110110011100111001110011111111111111111111111111"),
                ("1011010110101101011010110101101001110011010011101011010110101101001001110101101001001010010100101001100111001110011100111001111010110101101010011100111011010110101101011010110101101011010110101101011010110110011100111001110011111111111111111111111111"),
                ("1011010110101101011010110101101011010110100111001110011100111001110011100111001110011100111001110011100111001110011100111001111010110101101010011100111011010110101101011010011100111001110110101101011010110011001111011110111111111111111111111111111111"),
                ("1001110011100111001110011100111100111001101101011010110110011100101100110011100110011101101011010011101101011010011101101011010011100111101011001110011011010011100111100111001110011100110011100110110001100011001111111111111111111111111111111111111111"),
                ("1001110011100111001110011100111100111001101101011010110110011100101100110011100110011101101011010011101101011010011101101011010011100111101011001110011011010011100111100111001110011100110011100110110001100011001111111111111111111111111111111111111111"),
                ("1100111001110011100111001110011100111001100111100111001110011100101110111011110111001110011100111001110011100101100110011100110011100111100110011100111001111001110011100101100011001110101100011000110001100111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001110011100111001110011111011110111101111011110011100111011101011000110001100011100111001110011000110011001110011100111001110011001111001110010110001100011000111011110111101111111111111111111111111111111111111111111111111111111"),
                ("1100111001110011100111001110011100111001110011111011110111101111011110011100111011101011000110001100011100111001110011000110011001110011100111001110011001111001110010110001100011000111011110111101111111111111111111111111111111111111111111111111111111"),
                ("0111001110011001100111001110010110001100111101111011110111101111011111111111111111110011100111011110111101111011110111101111011001110011100111001110011100101100011001111011110111101111011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_2_2
                ("1111111111011101100111001110011001110011101101011010110100111001101001010000100001000010000100011011101111011100001101111011111011110111101101000010000100111000110001100001001010011101010110101101001110011110011111011110011001100111001011001111111111"),
                ("1111111111011101100111001110011001110011101101011010110100111001101001010000100001000010000100011011101111011100001101111011111011110111101101000010000100111000110001100001001010011101010110101101001110011110011111011110011001100111001011001111111111"),
                ("1111111111011001100111001110011001110011101101011010110110101101011010010010100101000110111101110111000010000100001000010000110111101111011101000010000100111000110000100101001010011101010011100111101011010100111100111001110011111011110011101111111111"),
                ("1111111111110011100111001110011001110011101101011010110100111001110011100111001101000101111011100001101111011110111101111011110111101111101101000010000100001000010001100001001010011101010110101101001110011110011111011110011001110111101111111111111111"),
                ("1111111111110011100111001110011001110011101101011010110100111001110011100111001101000101111011100001101111011110111101111011110111101111101101000010000100001000010001100001001010011101010110101101001110011110011111011110011001110111101111111111111111"),
                ("1111111111110011100111001110011001110011101101011010110110001100001001110001100001001010000100010111000010000100001000010000110111101111101101000010000100001000010000100101001010011101010011100111101011010100111100111001110011100111001111111111111111"),
                ("1111111111011001100111001110011100111001101101001110011100111001111010110001100001000110111101100001101111011101000101111011110111101111011101000010000100001000010000100101001010010100110011100111011010110101101011010110110011100111001110011111111111"),
                ("1111111111011001100111001110011100111001101101001110011100111001111010110001100001000110111101100001101111011101000101111011110111101111011101000010000100001000010000100101001010010100110011100111011010110101101011010110110011100111001110011111111111"),
                ("1111111111111101100111001100111011010110100110100101001100111001110011100111001101000101111011100001101111011110111000010000110111101111101101000010000100001000010000100101001010010100110011100111011010110101101100111001011001111011110111101111111111"),
                ("1111111111111101111011110110011011010110100111101011010110101101001001110001100001001010000100000001000010000100001101111011111011110111011101000010000100001000010000100001001010011100010011100111011010110101101001110011110010110001100111101111111111"),
                ("1111111111111101111011110110011011010110100111101011010110101101001001110001100001001010000100000001000010000100001101111011111011110111011101000010000100001000010000100001001010011100010011100111011010110101101001110011110010110001100111101111111111"),
                ("1111111111111101111011110110011100111001100111101011010110101101011000110101101001001010000100010111000010000100001110111101101000010000100001000010000100001000010000100001000010000100111010110101001110011101101011010110110011110111101111101111111111"),
                ("1111111111111101111011110110011100111001100111101011010110101101011000110101101001001010000100010111000010000100001110111101101000010000100001000010000100001000010000100001000010000100111010110101001110011101101011010110110011110111101111101111111111"),
                ("1111111111111111111011110011100110001100100110100101001110001100001000010010100101001010000100001000110111101111011010000100001000010000100001000010000100001000010000100001001010011001111010110101001110011101101100111001011001111011110111111111111111"),
                ("1111111111111110111001110111011100111001100111101011010010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110001011010110101101011010110101101100111001011001111111111111111111111111"),
                ("1111111111111110111001110111011100111001100111101011010010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100011000110001011010110101101011010110101101100111001011001111111111111111111111111"),
                ("1111111111111101110111101110011001110011100110100101001010000100001000010000100001000010000100001000010000100001000110111101110111101110100001000010000100001000010000100111010110101101011010110101101011010110101100111001011001111111111111111111111111"),
                ("1111111111011100110001100110011011010110100110100101001010000100001000010010100111000010010100101000010000100001000101111011100001000010100001000010000100001000010000100011010110101001111010110100100101001010011001110011011001111011110111111111111111"),
                ("1111111111011100110001100110011011010110100110100101001010000100001000010010100111000010010100101000010000100001000101111011100001000010100001000010000100001000010000100011010110101001111010110100100101001010011001110011011001111011110111111111111111"),
                ("1111111111111100110001100110011001110011100110100101001010010100111000010010100101001010000100011011110111101101000101111011100001000010100001000010000100001000010000100111010110101001110011100111001110011100111001110011110011110111101111011111111111"),
                ("1111111111111100111001110110011011010110100111001110011100111001111010010010100101000010000100010111000010000110111101111011111011110110100001000010000100101001010010100001001010010100111010110101011010110101101011010110101101100111001110011111111111"),
                ("1111111111111100111001110110011011010110100111001110011100111001111010010010100101000010000100010111000010000110111101111011111011110110100001000010000100101001010010100001001010010100111010110101011010110101101011010110101101100111001110011111111111"),
                ("1111111111111100111001110011001001110011100111001110011100111001111010010010100101001010000100010111000010000110111010000100001000010000100001000010001100001000010000100001001010010100111010110101001110011100111100111001100111100111001110011111111111"),
                ("1111111111111100110001100110011011010110100111001110011101101011010011010000100001000010000100001000101111011100001101111011101000010000100001000010000100101001010010100111000110001101010011100111001110011110011100111001110011100111001011001111111111"),
                ("1111111111111100110001100110011011010110100111001110011101101011010011010000100001000010000100001000101111011100001101111011101000010000100001000010000100101001010010100111000110001101010011100111001110011110011100111001110011100111001011001111111111"),
                ("1111111111110011100111001100111001110011110101101011010100111001101001010000100001000010010100101000010000100010111010000100001000010000100001001010011100011000110000100111010110101011010110101101100111001110011100111001110011100111001111111111111111"),
                ("1111111111110011100111001100111001110011110101101011010100111001101001010000100001000010010100101000010000100010111010000100001000010000100001001010011100011000110000100111010110101011010110101101100111001110011100111001110011100111001111111111111111"),
                ("1111111111110011100111001110011101011010110101101011010110101101001001010000100001000010010100101001010000100001000010000100001001010010100001001010010100001001010011101010011100111001110011100111100111001110011100111001110011111111111111111111111111"),
                ("1111111111110011100111001100111100111001100111001110011110101101001001010010100101001010010100101000010000100001000010000100001000010000100101000010000100001001010011001110110101101001110011100111001110011110011001110011110011111111111111111111111111"),
                ("1111111111110011100111001100111100111001100111001110011110101101001001010010100101001010010100101000010000100001000010000100001000010000100101000010000100001001010011001110110101101001110011100111001110011110011001110011110011111111111111111111111111"),
                ("1111111111110011001110011100111011010110101101011010110110101101001001110001100001000010000100001000010000100001000010000100001000010000100001001010010100001001010011001110110101101011010110101101011010110100111001110011110011111111111111111111111111"),
                ("1111111111011001100111001110011001110011101101011010110110101101001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010001001110110101101011010110101101011010110101101100111001110011111111111111111111111111"),
                ("1111111111011001100111001110011001110011101101011010110110101101001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010001001110110101101011010110101101011010110101101100111001110011111111111111111111111111"),
                ("1111111111111100110001100110011100111001101101011010110101101011010011110101101001000010000100001000010000100001001010010100101000010000100001000010000100101001010011011010110101101011010011100111001110011101101100111001011001111111111111111111111111"),
                ("1111111111111100110001100011001100111001100111011010110101101011010011110001100001000010000100001000010010100101001110001100001001010010100101001010010100110011100111011010110101101011011001110010110001100110011100111001111111111111111111111111111111"),
                ("1111111111111100110001100011001100111001100111011010110101101011010011110001100001000010000100001000010010100101001110001100001001010010100101001010010100110011100111011010110101101011011001110010110001100110011100111001111111111111111111111111111111"),
                ("1111111111111100111001110111011100111001100111011010110101101011010110110101101001001010000100001000010010100101001010010100111000110001101011000110000100111010110101001110011100111011001100011001111011110011001110111101111111111111111111111111111111"),
                ("1111111111111111111011110011001001110011101101011010110101101011010110101101011011000010000100001000010010100111000110001100011010110101011010011100111101010110101101011011001110011001111001110010110001100110010110001100111101111111111111111111111111"),
                ("1111111111111111111011110011001001110011101101011010110101101011010110101101011011000010000100001000010010100111000110001100011010110101011010011100111101010110101101011011001110011001111001110010110001100110010110001100111101111111111111111111111111"),
                ("1111111111111111111111111011000110001100101101011010110101101011010110100111001111000010000100001000110001100010011100111001110011100111011010011100111011010110101101011011001110011100111001110010111001110011001100111001100111111111111111111111111111"),
                ("1111111111111111111111111011000110001100101101011010110101101011010110100111001111000010000100001000110001100010011100111001110011100111011010011100111011010110101101011011001110011100111001110010111001110011001100111001100111111111111111111111111111"),
                ("1111111111111111111111111111110110001100011001100111001110011100111001101101011010110100111001111000100111001110110101101011010011100111001110011100111011010110101101011011001110011100111110111100111001110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111101100111001110011100111001110011100110011101101011010011100111001110110101101011010110101101011010110101101011010110101101001111001110011111011110111101111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111101100111001110011100111001110011100110011101101011010011100111001110110101101011010110101101011010110101101011010110101101001111001110011111011110111101111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111100111001011000110001100110011100110011101101011010110101101011010110100111001111001110011100111001110011100110011100111100101100011001111011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111101111011110110011100111001110011100110011101101011010110100111001111001110011100111001110010110001100011000110001110011101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111101111011110110011100111001110011100110011101101011010110100111001111001110011100111001110010110001100011000110001110011101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111101100011000110011001101101011010110100111001111001110011100111001110010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111001100110001100001100011000110011110111101100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111001100110001100001100011000110011110111101100111001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_2_3
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111110111101111011110011000110011001110011100111001110011100111110111101111011110111101111001110011101111011111111111111111110111101111011110111100110001100110011100111001011000111001110"),
                ("1111111111111111111111111111111111111111111111111111111111101111001110011000110001100110011100110011110011100111001110011100101100011000111001110011100110001100011001110101110011101111011110111101111011110110011100111001110011100111001110011100111001"),
                ("1111111111111111111111111111111111111111111111111111111111101111001110011000110001100110011100110011110011100111001110011100101100011000111001110011100110001100011001110101110011101111011110111101111011110110011100111001110011100111001110011100111001"),
                ("1111111111111111111111111111111111111111111110110001100011000110011101011000110011001110011100110011100111001111001100111001111001110010110011001110011100111001110011100111101111010111011001110011100111001100111100111001110011100111001110011100111001"),
                ("1111111111111111111111111111111111111111011000110001100100111001111001110011100111001100111001110110110011100111010100111001110110101101001110110101101001110110101101001111001110010110011001110011011010110101101100111001100111001110011100111001110011"),
                ("1111111111111111111111111111111111111111011000110001100100111001111001110011100111001100111001110110110011100111010100111001110110101101001110110101101001110110101101001111001110010110011001110011011010110101101100111001100111001110011100111001110011"),
                ("1111111111111111111111111111111111011110011001011010110101101011010011100111001110110101101011010110100111001111010110101101010011100111001110011100111001110011100111001110011100111001110011100111001110011100111011010110101101011010110101101011010110"),
                ("1111111111111111111111111110011100111001110011011010110101101011010110101101011010110101101011010110100111001111010110101101010011100111001110011100110100101001010010100111010110100100111010110101101011010010011001110011101101011010110101101011010110"),
                ("1111111111111111111111111110011100111001110011011010110101101011010110101101011010110101101011010110100111001111010110101101010011100111001110011100110100101001010010100111010110100100111010110101101011010010011001110011101101011010110101101011010110"),
                ("1111111111111111111011110011001100111001110011011010110101101011010110101101011010110110101101011010110101101011010100111001110110101101001110011100110100101000010000100001001010011100011010110101101011010100111001110011110001001110011110101001110011"),
                ("1111111111111111111011110011001100111001110011011010110101101011010110101101011010110110101101011010110101101011010100111001110110101101001110011100110100101000010000100001001010011100011010110101101011010100111001110011110001001110011110101001110011"),
                ("1111111111111111111011110011001100111001110011011010110101101011010110100111001110011010010100101001010010100101001010010100110011100111101011010110101100001000010000100001000010000100011000110000100101001100111101011010010011001110011110100100101001"),
                ("1111111111111111100111001110011100111001101101001110011101101011011010110001100011010010010100111000010010100101000010000100001000010000100101001010010100101001010010100001000010000100111010110101100011000100111100011000110001001110011010010100001000"),
                ("1111111111111111100111001110011100111001101101001110011101101011011010110001100011010010010100111000010010100101000010000100001000010000100101001010010100101001010010100001000010000100111010110101100011000100111100011000110001001110011010010100001000"),
                ("1111111111011001100111001100111001110011101101100011000110001100001001010000100001000010000100001000010010100101000010000100001000010000100101000010000100111000110000100001000010000100101001010010100101001010000100001000010010100001000010000100001000"),
                ("1111011110011001100111001101101011010110100110100001000010000100001000010000100001000010000100001000010010100101001010010100101000010000100001000010000100001001010010100001000010000100001000010000100001000101111101111011010001011110111110110100001000"),
                ("1111011110011001100111001101101011010110100110100001000010000100001000010000100001000010000100001000010010100101001010010100101000010000100001000010000100001001010010100001000010000100001000010000100001000101111101111011010001011110111110110100001000"),
                ("0110001100110011001110011101101001110011110000100001000010000100001000010000100001000010000100001000010000100001001010000100001000010001011110111101111101101000010000100001000010000100010111101110000100001000010000100001101110000100001101111101111011"),
                ("1100011000101101011010110101101001110011100111100011000010010100101001010010100101000010000100001000010000100001000010000100010111101110000100001000011101101000010000100001000010001101100001000010000100001101111011110111000011011110111000011011110111"),
                ("1100011000101101011010110101101001110011100111100011000010010100101001010010100101000010000100001000010000100001000010000100010111101110000100001000011101101000010000100001000010001101100001000010000100001101111011110111000011011110111000011011110111"),
                ("0110001100101101011010110101101011010110101101001110011110001100001001010010100101001010000100001000010000100001000101111011100001000011011110111101110100001000010000100001000010001101100001000010000100001101110100001000000011011110111000010000100001"),
                ("0110001100100111001110011100111011010110101101001110011110001100001001110001100001001010000100001000010000100001000010000100010111101110100010111101111011110111101111101101000010000100011011110111011110111000011011110111000011011110111000011011110111"),
                ("0110001100100111001110011100111011010110101101001110011110001100001001110001100001001010000100001000010000100001000010000100010111101110100010111101111011110111101111101101000010000100011011110111011110111000011011110111000011011110111000011011110111"),
                ("1111011110110011100111001110011011010110100111001110011110101101011000010010100101000010000100001000010000100001001010000100001000010000100011011110110000100001000011011101000010000100001000010001101111011101111011110111101111011110111101111101111011"),
                ("1111011110110011100111001110011011010110100111001110011110101101011000010010100101000010000100001000010000100001001010000100001000010000100011011110110000100001000011011101000010000100001000010001101111011101111011110111101111011110111101111101111011"),
                ("1100111001110011100111001110011011010110100111011010110101101011011010010010100101000010000100001000010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010001011110111110111011110111110111101111011101111101111011"),
                ("1100111001110011100111001110011011010110100111001110011100111001111000010010100101000010000100001001010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("1100111001110011100111001110011011010110100111001110011100111001111000010010100101000010000100001001010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000"),
                ("1111111111011000110001100110011011010110101101011010110110101101001001010010100101001010000100001000010000100001000110001100001001010011100001001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000010010100101001"),
                ("1111111111111110110001100100111011010110101101011010110101101011011010100111001101001010000100001001010010100101001110001100001001010010100001001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011000"),
                ("1111111111111110110001100100111011010110101101011010110101101011011010100111001101001010000100001001010010100101001110001100001001010010100001001010010100001000010000100001000010000100001000010000100001000010000100001000010000100001000110001100011000"),
                ("1111111111111110110001100110011001110011101101011010110101101011010011101101011010110100111001110011100111001111010010010100101001010010100001000010000100101000010000100101000010000100001000010000100001000010010100101001010011100011000010011100011000"),
                ("1111111111111110111001110011001100111001110011100111001110011100110011101101011010110101101011010110101101011010011110101101011000110000100101001010011101011010110101101011000110000100101000010000100101001010010100101001010010100101001010010100101001"),
                ("1111111111111110111001110011001100111001110011100111001110011100110011101101011010110101101011010110101101011010011110101101011000110000100101001010011101011010110101101011000110000100101000010000100101001010010100101001010010100101001010010100101001"),
                ("1111111111111111111111111111101111011110110011100111001100111001110110101101011010110101101011010110100111001110011101101011011010110100100101001010011001110011100111101010110101101001101001010011100011000010010100101001110101101011010110101101011010"),
                ("1111111111111111111111111111111111011110111101100111001110011100101100110011100110011101101011010110100111001110011101101011010011100111101011010110101001111010110101101010110101101101011010110101001110011100111001110011100111011010110100111011010110"),
                ("1111111111111111111111111111111111011110111101100111001110011100101100110011100110011101101011010110100111001110011101101011010011100111101011010110101001111010110101101010110101101101011010110101001110011100111001110011100111011010110100111011010110"),
                ("1111111111111111111111111111111111111111011100111001110011000110011110011000110010011101101011010110100111001111001110011100110011100111001110110101101001101001010011101010110101101001110011100111011010110101101011010110110101001110011110101001110011"),
                ("1111111111111111111111111111111111111111011100111001110011000110011110011000110010011101101011010110100111001111001110011100110011100111001110110101101001101001010011101010110101101001110011100111011010110101101011010110110101001110011110101001110011"),
                ("1111111111111111111111111111111111111111111110110001100110011100101100110011100110110101101011010011110011100111001110011100111001110011001110110101101001101001010011101010110101101011010110101101011010110101101011010110100111100111001100111100111001"),
                ("1111111111111111111111111111111111111111111111100111001011000110011101110011100111001110011100110011100111001111001110011100111001110011100110110101101001110011100111100111001110011100110110101101001110011110011011010110110011111011110110011111011110"),
                ("1111111111111111111111111111111111111111111111100111001011000110011101110011100111001110011100110011100111001111001110011100111001110011100110110101101001110011100111100111001110011100110110101101001110011110011011010110110011111011110110011111011110"),
                ("1111111111111111111111111111111111111111111111001110011111101111011111111111111101100110011100111001110011100111001110011100111001110011001110110101101100101100011000110001100011000110011001110011100111001011001100111001110010110001100110010110001100"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011110111110111101111111111111111111011101111010110001100111101100111001110011110111101111101100111001"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100111001110011100111001110011110111110111101111111111111111111011101111010110001100111101100111001110011110111101111101100111001"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011001100111001110011110111111111111111111111111111111111110111101111011110111101100111001111111111111111011100110001100"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_3_0
                ("1100111001111111111111111111111111111111111111111111111111111111111111111011110111001110011100111001110011100110011100111001110011100111100110011100110100101001010010100111010110101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1100111001111111111111111111111111111111111111111111111111111111111111111011110111001110011100111001110011100110011100111001110011100111100110011100110100101001010010100111010110101111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111110011100111001100111001110011100111001110110101101011010110101101100110011100111001110011100111101001100011001111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111011010110101101011011001110011100110110101101011010110101101011010110101101011010110101101011010011100111100111001110011100101100011000110011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111011010110101101011011001110011100110110101101011010110101101011010110101101011010110101101011010011100111100111001110011100101100011000110011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111101101011010110101101011010110100111001110011101101011010110101101011010110101101011010110101101011010011100111001110011100111011010011100111001110011100111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111011010110101101011010110100111001111010010010100111010101101011010110100111001110011101101011010011100111011010110101101001110110101101101011010110101011001100011001111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111011010110101101011010110100111001111010010010100111010101101011010110100111001110011101101011010011100111011010110101101001110110101101101011010110101011001100011001111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111001110011110101001110011100111001101001010010100111010100111001110110100111001110011101101011011010110101101011010110101001110110101101001111000110001001110110101100110001100011001111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111101011010010011101011010110101101001001110001100001001110001100001001100111001110110100111001111000110000100111000110001011010110101101101001001010011101010110101101100111001110010111001110111111111111111111111111111111"),
                ("1111111111111111111111111111111101011010010011101011010110101101001001110001100001001110001100001001100111001110110100111001111000110000100111000110001011010110101101101001001010011101010110101101100111001110010111001110111111111111111111111111111111"),
                ("1111111111111111111111111101101101011010010011100011000010000100001000010000100001000010010100101001110001100010011110001100001001010010100101001010011001110110101101101001001010011100010011100111001110011011001111011110101101111111111111111111111111"),
                ("1111111111111111111111111101101101011010010011100011000010000100001000010000100001000010010100101001110001100010011110001100001001010010100101001010011001110110101101101001001010011100010011100111001110011011001111011110101101111111111111111111111111"),
                ("1111111111111111100111001101101101011010010011100011000010010100101000010000100001000010000100001001110001100011010010010100101001010010100001000010000100001001010010100101001010011100001001010011101011010110011011010110101100110001100111111111111111"),
                ("1111111111111111001110011100111100011000010010100101001010010100101000010010100101001010000100001000010010100101001010010100101000010000100001000010000100001000010000100001001010010100101001010011001110011101101011010110101101100111001111111111111111"),
                ("1111111111111111001110011100111100011000010010100101001010010100101000010010100101001010000100001000010010100101001010010100101000010000100001000010000100001000010000100001001010010100101001010011001110011101101011010110101101100111001111111111111111"),
                ("1111111111111110110001100110011101011010010010100101001010000100001000010010100101001010010100101000010000100001000010010100101000010000100001000010000100001000010000100101001010010100010011100111011010110100111100111001011000110001100111111111111111"),
                ("1111111111111111111011110110011001110011110100100101001010010100101000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100111010110101011010110101101100111001110010110001100111111111111111"),
                ("1111111111111111111011110110011001110011110100100101001010010100101000010000100001001010010100101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100111010110101011010110101101100111001110010110001100111111111111111"),
                ("1111111111111111110111101110011011010110110100100101001010000100001000010010100101001010000100001000010000100001000010000100001000010000100011011110110100001000010000100001000010000100111010110101011010110101101011010110101101100111001111111111111111"),
                ("1111111111111101111011110100111011010110110100100101001010010100101000010000100001000010000100001000010000100001000010000100001000010001101111011110110100001000010000100001000010000100011010110101011010110101101011010110101101100111001111011111111111"),
                ("1111111111111101111011110100111011010110110100100101001010010100101000010000100001000010000100001000010000100001000010000100001000010001101111011110110100001000010000100001000010000100011010110101011010110101101011010110101101100111001111011111111111"),
                ("1111011110011001110111101101101011010110100111100011000010010100101001010000100001000010000100010111101111011111011010000100001000010001011111011110110100001000010000100001000010000100001000010001100011000110101101011010100111001110011011000110001100"),
                ("1111011110110011100111001011001011010110101101011010110110101101001001010010100101000010000100010111000010000110111000010000100001000011011110111101110100001000010000100001000010000100001000010000100001000010010100101001110101101011010110011100111001"),
                ("1111011110110011100111001011001011010110101101011010110110101101001001010010100101000010000100010111000010000110111000010000100001000011011110111101110100001000010000100001000010000100001000010000100001000010010100101001110101101011010110011100111001"),
                ("1100111001110011100111001100111001110011101101011010110110101101001000010000100001000010000100010111000010000110111101111011110111101110000110111101110100001000010000100001000010000100001000010000100001000010010100101001110101001110011110011100111001"),
                ("1100111001110011100111001100111001110011101101011010110110101101001000010000100001000010000100010111000010000110111101111011110111101110000110111101110100001000010000100001000010000100001000010000100001000010010100101001110101001110011110011100111001"),
                ("1100111001011001111011110111101100111001110011011010110110101101001000010000100001000110111101100001101111011100001101111011111011110111101100001000011101101000010000100001000010000100001000010000100001000010011100011000100111001110011110011100111001"),
                ("1111111111011000111001110111100110001100110011011010110100111001101000010000100011011000010000100001101111011110111101111011100001000010100010111101111011101000010000100001001010010100001000010000100101001110101001110011011000110001100110011111111111"),
                ("1111111111011000111001110111100110001100110011011010110100111001101000010000100011011000010000100001101111011110111101111011100001000010100010111101111011101000010000100001001010010100001000010000100101001110101001110011011000110001100110011111111111"),
                ("1111111111111111111011110111100110001100100110100101001010010100101000010000100011011101111011110111010000100001000101111011100001000010000100001000011101101000010000100101001010010100101001010010100101001100111011010110111100111001110111111111111111"),
                ("1111111111111111111011110011001100111001010010100001000010000100001001110001100001000110111101101000110111101110111101111011100001000010000100001000011101101000010000100001000010000100001000010000100101001100111011010110011001111011110111111111111111"),
                ("1111111111111111111011110011001100111001010010100001000010000100001001110001100001000110111101101000110111101110111101111011100001000010000100001000011101101000010000100001000010000100001000010000100101001100111011010110011001111011110111111111111111"),
                ("1111111111111110111001110111011001110011110000100001000010000100001001010010100101000010000100010111101111011110111000010000100001000011011100001000011101101000010000100001000010000100001000010000100001000110001001110011100111111011110111101111111111"),
                ("1111111111111110110001100110011001110011010000100001000010000100001000010000100011011110111101110111000010000100001000010000110111101111011100001000010000110111101110100001000010000100001000010000100001000010011101011010101101100111001011000110001100"),
                ("1111111111111110110001100110011001110011010000100001000010000100001000010000100011011110111101110111000010000100001000010000110111101111011100001000010000110111101110100001000010000100001000010000100001000010011101011010101101100111001011000110001100"),
                ("1111111111111111011010110101101001110011010010100001000010000100001000010000100001000110111101100001000010000100001101111011111011110111101101000010000100010111101111011111011110110100001000010000100001000010001101011010101101001110011110011100111001"),
                ("1111111111111111011010110101101011010110110100100001000010000100001000010000100001000010000100010111101111011110111101111011100001000011011101000010001011100001000010000100001000011101101000010000100001000010001101011010101101001110011110011100111001"),
                ("1111111111111111011010110101101011010110110100100001000010000100001000010000100001000010000100010111101111011110111101111011100001000011011101000010001011100001000010000100001000011101101000010000100001000010001101011010101101001110011110011100111001"),
                ("0111001110011001011010110100111001110011110100100101001010000100001000010000100001001010000100011011101111011110111000010000100001000010000110111101111011100001000011101101000010000100001000010000100001000010001001110011100110110001100111101111011110"),
                ("0111001110011001011010110100111001110011110100100101001010000100001000010000100001001010000100011011101111011110111000010000100001000010000110111101111011100001000011101101000010000100001000010000100001000010001001110011100110110001100111101111011110"),
                ("0110001100111101001110011110101100011000010010100001000010010100101001010000100001001010000100010111000010000100001000010000100001000011011111011110111011101000010000100001000010000100001000010000100001000010011011010110110011111011110111101111111111"),
                ("1100111001011001100111001100110100101001110000100001000010010100101001010000100011000010010100110111101111011100001000010000100001000010000110111101111101101000010000100001000010000100001000010000100001000010001001110011110011111011110111111111111111"),
                ("1100111001011001100111001100110100101001110000100001000010010100101001010000100011000010010100110111101111011100001000010000100001000010000110111101111101101000010000100001000010000100001000010000100001000010001001110011110011111011110111111111111111"),
                ("1100111001110011100111001100111101011010100110100101001010000100001001110001100001001010000100011011010000100010111000010000100001000010000100001000010000111011110110100001000010000100001001010010100101001010011001110011011000111001110111111111111111"),
                ("1100111001110011001110011100111011010110100110100101001010000100001000010010100101000010000100001000010000100010111000010000100001000010000100001000011011101000010000100001000010000100001000010001101011010100111001110011011001111011110111111111111111"),
                ("1100111001110011001110011100111011010110100110100101001010000100001000010010100101000010000100001000010000100010111000010000100001000010000100001000011011101000010000100001000010000100001000010001101011010100111001110011011001111011110111111111111111"),
                ("1111111111110011001110011101101001110011110000100101001010000100001000010000100001000010000100001000010000100011011101111011100001000010000100001000010000110111101110100001000010000100001000010001101011010101101011010110011000111001110111111111111111"),
                ("1111111111111111101011010100111101011010010011101011010010000100001000010000100001000010000100001000010000100001000101111011110111101110000100001000011011101000010000100001000010000100001000010001001110011101101011010110011000111001110111111111111111"),
                ("1111111111111111101011010100111101011010010011101011010010000100001000010000100001000010000100001000010000100001000101111011110111101110000100001000011011101000010000100001000010000100001000010001001110011101101011010110011000111001110111111111111111"),

                -- 7_explosion_3_1
                ("1111111111111111100111001110011100111001011000111001110111111111111111111111111111111111111111111111111111111111001110011100111110111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001"),
                ("1111111111111111100111001110011100111001011000111001110111111111111111111111111111111111111111111111111111111111001110011100111110111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001"),
                ("1111111111110011100111001110010110001100111100110001100111111111111111111111111111111111111111111111011000110001100110011100111001110010110011110111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1101011010100111001110011110011100111001100111011010110101101011010110011000110001110111101111011110011100111011110110011100111001110011110111110111101110111110111100110010011100111100111111111111111111111111111111111111111111111111111111111111111111"),
                ("1101011010100111001110011110011100111001100111011010110101101011010110011000110001110111101111011110011100111011110110011100111001110011110111110111101110111110111100110010011100111100111111111111111111111111111111111111111111111111111111111111111111"),
                ("1001110011101101001110011100111001110011110101001110011101101011010110110011100111101011000110011110111101111011110100111001101100011001011010011100111100111001110011100110011100111011010110101101111111111111111111111111111111111111111111111111111111"),
                ("1101011010100111011010110110100100101001110001001110011101101011010011100111001110011110011100101100011000110011001100111001110110101101011010110101101011010011100111101011000110001101011010110101101011010100111011010110111111111111111111111111111111"),
                ("1101011010100111011010110110100100101001110001001110011101101011010011100111001110011110011100101100011000110011001100111001110110101101011010110101101011010011100111101011000110001101011010110101101011010100111011010110111111111111111111111111111111"),
                ("0100101001110001001110011100111100011000010011101011010110101101001001010000100011000010010100110011110011100111001101101011010110101101001111010110101101011010110100100101001010010100101001010010100101001110101011010110101101111111111111111111111111"),
                ("1101011010010010100101001010010100001000010000100101001010000100001000010000100001000010000100001001101101011010110101101011010110101101100001001010010100101001010010100101001010011100011000110001101011010100111011010110101101011010110111111111111111"),
                ("1101011010010010100101001010010100001000010000100101001010000100001000010000100001000010000100001001101101011010110101101011010110101101100001001010010100101001010010100101001010011100011000110001101011010100111011010110101101011010110111111111111111"),
                ("0100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001001100111001111010110101101011010110100100101001010010100001001010010100001001010010100101000010001101011010100111001110011101101011010110111111111111111"),
                ("0100001000010000100001000010000100101001010010100001000010000100001000010000100001000010000100001001100111001111010110101101011010110100100101001010010100001001010010100001001010010100101000010001101011010100111001110011101101011010110111111111111111"),
                ("0100001000010000100001000010010100101001010010100001000010000100001000010000100001001010010100101000010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100101001010011101011010101101100111001111111111111111"),
                ("0100001000010000100101001110000100001000010000100001000010000100001000010000100001001110001100001000010000100001000010000100001001010010100001000010000100101000010000100101001010010100001000010001100011000010010100101001100111100111001110011110111101"),
                ("0100001000010000100101001110000100001000010000100001000010000100001000010000100001001110001100001000010000100001000010000100001001010010100001000010000100101000010000100101001010010100001000010001100011000010010100101001100111100111001110011110111101"),
                ("0100001000010000100001000010011100011000010010100101001010000100001000110111101101000010000100011011110111101101000010000100001000010000100001000010000100101001010010100101001010010100001000010000100101001110101101011010100111011010110110011100111001"),
                ("0100001000010000100001000010000100101001010000100001000010000100011011110111101101000110111101110111000010000111011010000100001000010000100001000010000100001001010010100101000010000100001001010011100011000100111011010110101101011010110100111100111001"),
                ("0100001000010000100001000010000100101001010000100001000010000100011011110111101101000110111101110111000010000111011010000100001000010000100001000010000100001001010010100101000010000100001001010011100011000100111011010110101101011010110100111100111001"),
                ("0100001000010000100001000110111011110111101111101111011101111011100001101111011110111010000100010111000010000100001101111011110111101111011101000010000100001000010000100001000010000100101001010010100101001101101011010110101101011010110100111100111001"),
                ("0100001000010000100001000010001011110111000011011110111101111011100001000010000110111110111101101000101111011110111000010000100001000011011101000010000100001000010000100001001010011100011000110001001110011100111001110011101101011010110100111100111001"),
                ("0100001000010000100001000010001011110111000011011110111101111011100001000010000110111110111101101000101111011110111000010000100001000011011101000010000100001000010000100001001010011100011000110001001110011100111001110011101101011010110100111100111001"),
                ("0100001000110111011110111101110000100001000011011110111101111011100001000010000110111101111011101000101111011100001101111011110111101111101101000010000100001000010000100001001010011101010011100111011010110100111001110011101101011010110101101001110011"),
                ("1011110111101110000100001000010000100001000010000100001101111011110111000010000100001101111011110111101111011110111101111011100001000010100001000010000100001000010000100101001010010100111000110001001110011101101011010110101101011010110101101001110011"),
                ("1011110111101110000100001000010000100001000010000100001101111011110111000010000100001101111011110111101111011110111101111011100001000010100001000010000100001000010000100101001010010100111000110001001110011101101011010110101101011010110101101001110011"),
                ("1011110111000010000100001000010000100001000010000100001000010000111011101111011100001000010000100001000010000111011101111011100001000010100001000010000100001000010000100001000010000100101001010011100011000110101001110011101101011010110101101001110011"),
                ("1011110111000010000100001000010000100001000010000100001000010000111011101111011100001000010000100001000010000111011101111011100001000010100001000010000100001000010000100001000010000100101001010011100011000110101001110011101101011010110101101001110011"),
                ("0000100001000010000100001000010000100001101110000100001101111011111011101111011110111000010000100001010000100011011000010000110111101111011111011110110100001000010000100001000010000100001001010010100101001110101011010110101101011010110110011100111001"),
                ("0000100001000010000100001000011011110111110111011110111010000100001000000010000100001000010000100001101111011100001101111011110111101111101111011110111101101000010000100001000010000100001001010011100011000110101011010110100111001110011100111001110011"),
                ("0000100001000010000100001000011011110111110111011110111010000100001000000010000100001000010000100001101111011100001101111011110111101111101111011110111101101000010000100001000010000100001001010011100011000110101011010110100111001110011100111001110011"),
                ("1011110111000011011110111000011101111011101111011110111101111011101000000010000111011110111101111011101111011111011010000100001000010000100001000010000100001000010000100001000010000100010011100111011010110100111001110011100111100111001100110100101001"),
                ("0100001000101110100001000110110100001000010000000100001000010000110111101111011101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100110110101101011010110101101011010110100111100111001100110100101001"),
                ("0100001000101110100001000110110100001000010000000100001000010000110111101111011101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100110110101101011010110101101011010110100111100111001100110100101001"),
                ("0100001000010000100001000010000100001000010001101111011000010000110111010000100001000010000100001001010000100001000010000100001000010000100001000010000100001000010000100101000010000100111010110101101011010100111101011010101101100111001110100100101001"),
                ("0100001000010000100001000010000100001000010000100001000000010000111011010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100101001010010100101001010010100101001110001101011010100110110001100011001101011010"),
                ("0100001000010000100001000010000100001000010000100001000000010000111011010000100001000010000100001001010010100101000010000100001000010000100001000010000100001000010000100101001010010100101001010010100101001110001101011010100110110001100011001101011010"),
                ("0100001000010000100001000010000100001000010000100001000110111101101000010000100001000010000100001001010000100001000010000100001000010000100001000010000100101001010010100001001010011100011000110001101011010100111011010110100110110001100111111111111111"),
                ("0100001000010000100001000010010100001000010000100001000010000100001000010000100001000010000100001001010000100001000010000100001000010000100011010110101101011010110101001101001010010100110011100111011010110101100110001100100111111111111111111111111111"),
                ("0100001000010000100001000010010100001000010000100001000010000100001000010000100001000010000100001001010000100001000010000100001000010000100011010110101101011010110101001101001010010100110011100111011010110101100110001100100111111111111111111111111111"),
                ("1001110011110101101011010010010100001000010000100001000010000100001000010000100001000010010100101001010010100101000010000100001000010001100010110101101011010110101101011010011100111101010011100111100111001011001111011110111111111111111111111111111111"),
                ("1001110011110101101011010010010100001000010000100001000010000100001000010000100001000010010100101001010010100101000010000100001000010001100010110101101011010110101101011010011100111101010011100111100111001011001111011110111111111111111111111111111111"),
                ("1011010110101101001110011010010100001000010010100001000010000100001000010010100111000100111001110011110101101001001010010100101001010011101010110101101011010110101101001110110101101100101100011001100111001011001111111111111111111111111111111111111111"),
                ("1011010110101101001110011100111001110011101101001110011110101101011010110101101010011101101011010110100111001111000010010100101001010011101010110101101011011001110011100110110101101011011110111100111001110111111111111111111111111111111111111111111111"),
                ("1011010110101101001110011100111001110011101101001110011110101101011010110101101010011101101011010110100111001111000010010100101001010011101010110101101011011001110011100110110101101011011110111100111001110111111111111111111111111111111111111111111111"),
                ("0110001100011000110001100011001100111001110011001110011101101011010110101101011010011011000110011110011000110010011110101101011010110101001110110101101011011001110010110010110101101011010110101101111111111111111111111111111111111111111111111111111111"),
                ("0111001110011101111011110011101111011110111100110001100100111001110011110011100111110111101111001110011000110010011100111001111010110101001111001110011100101100011000110011001110010110011111111111111111111111111111111111111111111111111111111111111111"),
                ("0111001110011101111011110011101111011110111100110001100100111001110011110011100111110111101111001110011000110010011100111001111010110101001111001110011100101100011000110011001110010110011111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111101111011110110011100111001011000110011110111111111111111110011100111001110011100111001110010110011101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110110011100111001011000110011111111111111111111111111111111001110011100111001110010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110110011100111001011000110011111111111111111111111111111111001110011100111001110010110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),

                -- 7_explosion_3_2
                ("1111111111111110111001110011001011010110101101001110011010000100001000010000100001000010000100010111000010000100001101111011110111101110100001000010000100001000010000100001000010000100001000010001101011010010011101011010100111101011010111111111111111"),
                ("1111111111111110111001110011001011010110101101001110011010000100001000010000100001000010000100010111000010000100001101111011110111101110100001000010000100001000010000100001000010000100001000010001101011010010011101011010100111101011010111111111111111"),
                ("1111111111111110111001110011001011010110101101101011010010000100001000010000100001000101111011100001000010000100001000010000110111101111101101000010000100001000010000100001000010000100001000010000100101001110001001110011101101001110011110011111111111"),
                ("1111111111111111111011110011001001110011100111101011010010000100001000010000100001000010000100010111000010000100001000010000100001000011011101000010000100001000010000100001001010010100001000010000100101001100111011010110100111001110011110011100111001"),
                ("1111111111111111111011110011001001110011100111101011010010000100001000010000100001000010000100010111000010000100001000010000100001000011011101000010000100001000010000100001001010010100001000010000100101001100111011010110100111001110011110011100111001"),
                ("1111111111111110111001110011001001110011010010100101001010010100101000010000100001000110111101100001000010000100001000010000100001000011011101000010001101101000010000100111000110000100101000010000100101001100111101011010100111100111001110011100111001"),
                ("1111111111111111111011110110011001110011010000100001000010000100001000010000100001000010000100011011101111011100001000010000100001000010000110111101111011101001010011100001000010000100101001010010100001000110000100101001100111100111001011001100111001"),
                ("1111111111111111111011110110011001110011010000100001000010000100001000010000100001000010000100011011101111011100001000010000100001000010000110111101111011101001010011100001000010000100101001010010100001000110000100101001100111100111001011001100111001"),
                ("1111111111111101111011110110011011010110010010100001000010000100001000010000100001000010000100010111110111101110111000010000100001000010000100001000011011101000010000100101000010000100101001010010100001000010011100011000110101001110011111100110001100"),
                ("1111011110111100110001100100111001110011010000100001000010000100001000010000100011011000010000110111101111011100001000010000100001000011011110111101111101101000010000100101000010000100001000010000100101001110101001110011100111011010110011000111001110"),
                ("1111011110111100110001100100111001110011010000100001000010000100001000010000100011011000010000110111101111011100001000010000100001000011011110111101111101101000010000100101000010000100001000010000100101001110101001110011100111011010110011000111001110"),
                ("1100111001110011001110011101101101011010010000100001000010000100011011000010000100001000010000110111010000100010111000010000110111101111011110111101111011101000010000100001000010000100001000010000100001000110101011010110101101011010110111111111111111"),
                ("1100111001110011001110011101101101011010010000100001000010000100011011000010000100001000010000110111010000100010111000010000110111101111011110111101111011101000010000100001000010000100001000010000100001000110101011010110101101011010110111111111111111"),
                ("1100111001110011001110011101101101011010010000100001000010000100001000110111101110111101111011101000010000100011011110111101110111101110000100001000010000111011110110100001000010000100001000010000100001000010011001110011101101011010110111111111111111"),
                ("0110001100011001100111001101101101011010010010100001000010000100001000010000100001000101111011100001000010000110111101111011100001000010000100001000011011111011110111101101000010000100001000010000100001000010001001110011110010110001100111111111111111"),
                ("0110001100011001100111001101101101011010010010100001000010000100001000010000100001000101111011100001000010000110111101111011100001000010000100001000011011111011110111101101000010000100001000010000100001000010001001110011110010110001100111111111111111"),
                ("1111111111111101111011110100111001110011110000100001000010000100001000010000100001000010000100011011000010000110111000010000100001000011011110111101111011101000010000100001001010010100101000010000100001000110001001110011111010111001110111111111111111"),
                ("1111111111111111111011110011001011010110100110100101001010000100001000010000100001000010000100011011000010000100001000010000110111101111011111011110110100011011110110100011000110000100101000010000100001000010011100111001011001111011110111111111111111"),
                ("1111111111111111111011110011001011010110100110100101001010000100001000010000100001000010000100011011000010000100001000010000110111101111011111011110110100011011110110100011000110000100101000010000100001000010011100111001011001111011110111111111111111"),
                ("1111111111111110111001110111101011010110100110100101001010010100101001010010100101001010000100011011000010000100001000010000110111101110100001000010001011110111101111101101000010000100001001010010100101001100110110001100111101111011110111111111111111"),
                ("1111111111110010110001100011001001110011110100100101001010000100001000010010100101000010000100010111101111011101000000010000110111101111011110111101110000100001000011101101000010000100010011100111011010110110010110001100111100111001110011001111111111"),
                ("1111111111110010110001100011001001110011110100100101001010000100001000010010100101000010000100010111101111011101000000010000110111101111011110111101110000100001000011101101000010000100010011100111011010110110010110001100111100111001110011001111111111"),
                ("1100111001110011001110011100111100011000010010100001000010000100001000010000100001000010000100011011000010000111011110111101110111101110000110111101110000111011110110100001000010000100011010110101011010110110011100111001111101111011110011001100111001"),
                ("1100111001110011001110011110100100101001010010100001000010000100001000010000100001000010000100001000101111011100001101111011110111101111011100001000011011101000010000100001000010000100011010110101011010110101101001110011100111100111001110011100111001"),
                ("1100111001110011001110011110100100101001010010100001000010000100001000010000100001000010000100001000101111011100001101111011110111101111011100001000011011101000010000100001000010000100011010110101011010110101101001110011100111100111001110011100111001"),
                ("1100111001110011101011010110100100101001010010100001000010000100001000010000100001000010000100001000101111011110111000010000100001000011011100001000011011101000010000100001001010010100111010110101011010110101101011010110011001100111001110011111011110"),
                ("1100111001110011101011010110100100101001010010100001000010000100001000010000100001000010000100001000101111011110111000010000100001000011011100001000011011101000010000100001001010010100111010110101011010110101101011010110011001100111001110011111011110"),
                ("0110001100011001001110011100111101011010110101100011000010000100001000010000100001000010000100001000110111101110111010000100001000010001101110111101111011101000010000100001000010000100101001010011100011000100111011010110101101110111101011001111011110"),
                ("1111111111111011100111001101101011010110101101011010110110101101001000010000100001000010000100001000110111101111011010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001110101011010110100111111011110111101111111111"),
                ("1111111111111011100111001101101011010110101101011010110110101101001000010000100001000010000100001000110111101111011010000100001000010000100001000010000100001000010000100001000010000100001001010010100101001110101011010110100111111011110111101111111111"),
                ("1111111111111111100111001101101011010110101101011010110110101101001001010000100001000010000100001000110111101101000010000100001000010000100001000010000100001000010000100101001010010100001000010000100101001110101011010110110011110111101111111111111111"),
                ("1111111111111110110001100110011100111001101101011010110110101101001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100001001010010100101001110101001110011110011111011110111111111111111"),
                ("1111111111111110110001100110011100111001101101011010110110101101001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001001010010100101000010000100001001010010100101001110101001110011110011111011110111111111111111"),
                ("1111111111111110110001100011001100111001100111011010110100111001101000010010100101001010000100001000010000100001000010000100001001010010100001000010000100001001010010100101001010010100001000010000100101001010011101011010110010110001100111111111111111"),
                ("1111111111111111100111001101101011010110101101001110011010010100101001010010100101000010000100001000010000100001000010000100001001010010100101001010010100001000010000100101001010010100001001010010100101001010011100011000100111001110011111111111111111"),
                ("1111111111111111100111001101101011010110101101001110011010010100101001010010100101000010000100001000010000100001000010000100001001010010100101001010010100001000010000100101001010010100001001010010100101001010011100011000100111001110011111111111111111"),
                ("1111111111111110110001100101101011010110110011101011010010010100111000010010100101001010010100101000010000100001000010010100101001010011101011000110000100101000010000100001000010000100001001010011100011000010011101011010101101100111001111111111111111"),
                ("1111111111111111111111111101101111011110011001001110011100111001111000010010100111010101101011010011010010100101001010010100111000110001001111000110000100101001010010100001000010000100001000010001100011000010011101011010101101111111111111111111111111"),
                ("1111111111111111111111111101101111011110011001001110011100111001111000010010100111010101101011010011010010100101001010010100111000110001001111000110000100101001010010100001000010000100001000010001100011000010011101011010101101111111111111111111111111"),
                ("1111111111111111111111111111110111001110110011100111001101101011011010010010100111010101101011010110110001100001001110001100010011100111011010011100110100111000110000100111000110000100111010110101101011010010011101011010111111111111111111111111111111"),
                ("1111111111111111111111111111110111001110110011100111001101101011011010010010100111010101101011010110110001100001001110001100010011100111011010011100110100111000110000100111000110000100111010110101101011010010011101011010111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111011000110001100101101011010011110001100010011101101011010011110101101011010110101101010110101101001110011100111011010011100111101001001010010100110011100111001110011110101001110011111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110011000110010110110101101011010101101011010011101101011010110100111001110110101101001110011100111011010110101101101001001010011101010011100111011010110101101011010110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111011110011000110010110110101101011010101101011010011101101011010110100111001110110101101001110011100111011010110101101101001001010011101010011100111011010110101101011010110111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111100111001110011100111001110110100111001110011100111001110110101101011010110101101011010110101101011010110101101001110011100111011010110101101011010110101101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111101100011000110011001110011100111001100111001110110101101011010110101101011010110101101011010110101101011011001110011100110110101101011010110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111101100011000110011001110011100111001100111001110110101101011010110101101011010110101101011010110101101011011001110011100110110101101011010110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111011000110011010100111001110011100111001111001101101011010110101101011010011100111001110011100111100111001110011111111111111111111111111111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111110101101001001010010100101001100111001111001100111001110011100111001111001110011100111001110011100111101111011111111111111111111111111111111111111111111111111111111111111100111001"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111110101101001001010010100101001100111001111001100111001110011100111001111001110011100111001110011100111101111011111111111111111111111111111111111111111111111111111111111111100111001"),

                -- 7_explosion_3_3
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100110011100111001110011100111111111111111111111111111111101100011001100111001110011111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100110011100111001110011100111111111111111111111111111111101100011001100111001110011111011110111111111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110101100110011100111001110011100111001110011111111111111111111001100011001100111001110011111011110111101111111111111111111111111111111111111111"),
                ("1111111111111111111111111111111111111111111111111111111111111111101100110011100101100011000110011001110011100110011110101101010011100111001101100011000111011110111101111011001110011001110011100110110001100111101111011110011101111011110011100111001110"),
                ("1111111111111111111111111111111111111111111111111111111111111111101100110011100101100011000110011001110011100110011110101101010011100111001101100011000111011110111101111011001110011001110011100110110001100111101111011110011101111011110011100111001110"),
                ("1111111111111111111111111111111111111111111111111111111101101011010110101101011001100110011100110110101101011010011110101101011010110101001101100011001111001100011001001110110101101011010110101101001110011110011100111001011000110001100011000110001100"),
                ("1111111111111111111111111111111111111111111110111001110111101111010110101101011011001110011100110110101101011011010010010100101001010011100010011100111011010110101101001111010110101101011010110101001110011101101001110011100111001110011101101011010110"),
                ("1111111111111111111111111111111111111111111110111001110111101111010110101101011011001110011100110110101101011011010010010100101001010011100010011100111011010110101101001111010110101101011010110101001110011101101001110011100111001110011101101011010110"),
                ("1111111111111111111111111111111111111111011001100111001011000110011001101101011010011101101011010110101101011011010010010100101001010010100111010110101001110011100111100001001010010100001000010000100001000010010100001000010011001110011101101011010110"),
                ("1111111111111111111111111111111111011110011001100111001100111001111010100111001110110101101011010110101101011011000010000100001000010000100001001010010100101001010010100001000010000100001000010000100001000010000100001000010011101011010110101001110011"),
                ("1111111111111111111111111111111111011110011001100111001100111001111010100111001110110101101011010110101101011011000010000100001000010000100001001010010100101001010010100001000010000100001000010000100001000010000100001000010011101011010110101001110011"),
                ("1111111111111111111111111100110110001100101101011010110100111001101001010010100110011110101101011010110101101001000010000100001000010000100001000010000100101000010000100001000010000100001000010000100001000010000100001000010010100001000010000100001000"),
                ("1111111111111111111111111100110110001100101101011010110100111001101001010010100110011110101101011010110101101001000010000100001000010000100001000010000100101000010000100001000010000100001000010000100001000010000100001000010010100001000010000100001000"),
                ("1111111111111110110001100100111011010110100111101011010110001100011000010010100101000010010100101001010000100001000010000100001000010000100001000010000100101000010000100001000010000100011011110110100001000010000100001000010000100001000010000100001000"),
                ("1101011010011000110001100100111101011010110000100101001010010100101001010010100101001010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010001101100001000010100001000010000100001000010000100001000010000100001000"),
                ("1101011010011000110001100100111101011010110000100101001010010100101001010010100101001010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010001101100001000010100001000010000100001000010000100001000010000100001000"),
                ("0100101001110101100111001101101101011010100111101011010110101101001001010000100001001010000100001000010000100001000010000100001000010000100001000010000100101000010000100001000010001011100001000011101111011010000100001000010000100001000010000100001000"),
                ("0100101001100111100111001100111011010110101101011010110101101011001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100010111101111011100001000010000100001010000100001000110110100001000101110100001000"),
                ("0100101001100111100111001100111011010110101101011010110101101011001001010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100010111101111011100001000010000100001010000100001000110110100001000101110100001000"),
                ("0100101001100111100111001100111001110011100111011010110100111001101000010000100001000010000100001000010000100001000010000100001000010001101110111101111101111011110111101100001000010100010111101111011110111101111101111011000011011110111000011011110111"),
                ("1001110011100111001110011100111011010110110101100011000010010100101000010000100001000010000100011011110111101111011101111011110111101110000110111101110000100001000010000100001000010100001000010001011110111110111011110111000010000100001000010000100001"),
                ("1001110011100111001110011100111011010110110101100011000010010100101000010000100001000010000100011011110111101111011101111011110111101110000110111101110000100001000010000100001000010100001000010001011110111110111011110111000010000100001000010000100001"),
                ("1100111001110011011010110101101011010110110100100101001010010100101000010000100001000010000100001000110111101110111101111011100001000011101101000010000000100001000011011110111101111101110111101110000100001101110000100001000010000100001000010000100001"),
                ("1001110011101101011010110101101001110011110101100011000010010100101001010000100001000010000100001000010000100001000000010000110111101111101100001000010000100001000010000110111101111101100001000010000100001000010000100001000010000100001000011011110111"),
                ("1001110011101101011010110101101001110011110101100011000010010100101001010000100001000010000100001000010000100001000000010000110111101111101100001000010000100001000010000110111101111101100001000010000100001000010000100001000010000100001000011011110111"),
                ("1001110011101101011010110101101011010110101101001110011110001100001001010010100101001010000100001000010000100001000000010000110111101111011110111101111011110111101110000100001000011011110111101110000100001000010000100001000010000100001101111011110111"),
                ("1001110011101101011010110101101011010110101101001110011110001100001001010010100101001010000100001000010000100001000000010000110111101111011110111101111011110111101110000100001000011011110111101110000100001000010000100001000010000100001101111011110111"),
                ("1001110011101101011010110101101001110011100111011010110100111001111010010010100101000010000100001000010000100011011101111011110111101110000110111101110100010111101111011100001000010000110111101111011110111000010000100001101111011110111110110100001000"),
                ("1100111001100111011010110101101001110011100111001110011110001100011000010010100101000010000100001000010000100010111000010000100001000011011110111101110100011011110111011100001000010000110111101111011110111000011011110111010000100001000010000100001000"),
                ("1100111001100111011010110101101001110011100111001110011110001100011000010010100101000010000100001000010000100010111000010000100001000011011110111101110100011011110111011100001000010000110111101111011110111000011011110111010000100001000010000100001000"),
                ("1100111001100111011010110101101011010110101100100101001010010100101001010000100001000010000100001000010000100010111101111011110111101110000100001000011011101000010001011110111101110000110111101111101111011101111011110111110110100001000010000100001000"),
                ("1100111001100111011010110101101011010110100111100011000010010100101000010000100001001010010100101000010000100001000010000100001000010001101100001000011011111011110110100011011110111101101000010000100001000010000100101001010000100001000010000100001000"),
                ("1100111001100111011010110101101011010110100111100011000010010100101000010000100001001010010100101000010000100001000010000100001000010001101100001000011011111011110110100011011110111101101000010000100001000010000100101001010000100001000010000100001000"),
                ("1100111001110011011010110100111101011010110100100101001010000100001000010010100101001010010100101001010000100001000010000100001000010000100011011110111101101000010000100011011110110100001000010000100101001010011100011000010010100001000010000100001000"),
                ("1110111101110011100111001100110100101001010011100011000010000100001000010010100101001010000100001001010000100001000010010100101000010000100001000010000100011000110000100101000010000100001000010000100001000010000100001000110000100101001010000100001000"),
                ("1110111101110011100111001100110100101001010011100011000010000100001000010010100101001010000100001001010000100001000010010100101000010000100001000010000100011000110000100101000010000100001000010000100001000010000100001000110000100101001010000100001000"),
                ("1111111111111111100111001101101101011010010010100101001010000100001000010000100001000010000100001000010000100001001010010100101000010000100001000010000100001001010010100101000010000100001000010000100001000010010100101001010010100001000010000100001000"),
                ("1111111111111111011010110101101001110011100111101011010010000100001001010010100101000010010100101000010010100101001110101101011010110101101010011100110100101000010000100001000010000100001000010000100001000010010100101001010000100001000010000100001000"),
                ("1111111111111111011010110101101001110011100111101011010010000100001001010010100101000010010100101000010010100101001110101101011010110101101010011100110100101000010000100001000010000100001000010000100001000010010100101001010000100001000010000100001000"),
                ("1111111111111111011010110101101011010110100111101011010110001100011000010010100101001010010100101001010010100111000101101011010110101101011010110101100100101000010000100001000010000100001000010000100101001010000100001000010010100101001010011101011010"),
                ("1111111111111111011010110101101011010110100111101011010110001100011000010010100101001010010100101001010010100111000101101011010110101101011010110101100100101000010000100001000010000100001000010000100101001010000100001000010010100101001010011101011010"),
                ("1111111111111111111111111101101011010110110100100101001010010100101001010010100101001110101101011010110101101010011101101011010110101101100111001110011001101001010011100001000010000100111010110101101011010010011100011000100111001110011110000100101001"),
                ("1111111111111111111111111111111011010110100111101011010110101101011010110001100011010100111001110110101101011010110101101011010011100111100101100011000110011001110011001110011100111001110110101101001110011110000100101001110101011010110100111101011010"),
                ("1111111111111111111111111111111011010110100111101011010110101101011010110001100011010100111001110110101101011010110101101011010011100111100101100011000110011001110011001110011100111001110110101101001110011110000100101001110101011010110100111101011010"),
                ("1111111111111111111111111111111111111111111111111111111101101011010110100111001111001110011100111001100111001110110011000110010011100111111011110111101111001100011001110111001110011011010110101101001110011110101001110011100111001110011101101001110011"),
                ("1111111111111111111111111111111111111111111111111111111111111111111001100111001101100111101111011101111101111011101110011100111001110011111001110011101111011110111100111001100011001011010110101101011010110100111100111001110011001110011100111101011010"),
                ("1111111111111111111111111111111111111111111111111111111111111111111001100111001101100111101111011101111101111011101110011100111001110011111001110011101111011110111100111001100011001011010110101101011010110100111100111001110011001110011100111101011010"),
                ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111001100110011100111001110010110001100011001111111111111111111111111111111111111111111110110001100111100110001100110011100111001110011111111111"),
                ("1100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111011001110011100111111111111111111111111111111111111111111111111111111110111001110011001100111001110011100111001111111111111111"),
                ("1100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111011001110011100111111111111111111111111111111111111111111111111111111110111001110011001100111001110011100111001111111111111111"),

                -- 8_bonus-life
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110001101011010110101101011010110111100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110001101011010110101101011010110111100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110001101011010110101101011010110111100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101101001010010100100111001110011110001100011000110001100010011100111001110100101001010010100101001010010011100111001101001010011101011010110101001110011100111010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101101001010010100100111001110011110001100011000110001100010011100111001110100101001010010100101001010010011100111001101001010011101011010110101001110011100111010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101101001010010100100111001110011110001100011000110001100010011100111001110100101001010010100101001010010011100111001101001010011101011010110101001110011100111010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011100111001110011010010100100111001110011010010100101001010000100001000010000100001001010010100110011100111001110011100111001101001010010100101000010001111011110111101101011010110101001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100100111001110011010010100101001010000100001000010000100001001010010100110011100111001110011100111001101001010010100101000010001111011110111101101011010110101001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100100111001110011010010100101001010000100001000010000100001001010010100110011100111001110011100111001101001010010100101000010001111011110111101101011010110101001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001000010000100001000010000100001010000100001000010000100011010110101101011000110001100001000010000100001110011100101101011010111111011110111101101011010110101010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001000010000100001000010000100001010000100001000010000100011010110101101011000110001100001000010000100001110011100101101011010111111011110111101101011010110101010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001000010000100001000010000100001010000100010100101001010011101111011110110100101001010011101111011110100100001000111001110011100100001000010000100101001010011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001000010000100001000010000100001010000100010100101001010011101111011110110100101001010011101111011110100100001000111001110011100100001000010000100101001010011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001000010000100001000010000100001010000100010100101001010011101111011110110100101001010011101111011110100100001000111001110011100100001000010000100101001010011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001010000100001000010000100001000101001010010100101001010000100001000010010000100001000000000000000000011101111010100001000010000100001000010000100101001010011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001010000100001000010000100001000101001010010100101001010000100001000010010000100001000000000000000000011101111010100001000010000100001000010000100101001010011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010010100101001010000100001000010000100001000101001010010100101001010000100001000010010000100001000000000000000000011101111010100001000010000100001000010000100101001010011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100100111001110011010000100001000101111011110111101001010000111001110011100101001010010101111011110111111101111011110110100101000100001000010000100001000010001001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100100111001110011010000100001000101111011110111101001010000111001110011100101001010010101111011110111111101111011110110100101000100001000010000100001000010001001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100100111001110011010000100001000101111011110111101001010000111001110011100101001010010101111011110111111101111011110110100101000100001000010000100001000010001001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101101001010010100010010100101001010000100001000111001110000110001100011001111011110111101110011100111011101111011110111100111000100001000010000100101001010011010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101101001010010100010010100101001010000100001000111001110000110001100011001111011110111101110011100111011101111011110111100111000100001000010000100101001010011010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101101001010010100010010100101001010000100001000111001110000110001100011001111011110111101110011100111011101111011110111100111000100001000010000100101001010011010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100100111001110011110001100011000101001010000000000000000011101111011110111101111011110111100111001110010100101001100011000110001001110011100111110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100100111001110011110001100011000101001010000000000000000011101111011110111101111011110111100111001110010100101001100011000110001001110011100111110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100100111001110011110101101010100101001010011100111001110011100111001110010100101001010011010110101001110011100111010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100100111001110011110101101010100101001010011100111001110011100111001110010100101001010011010110101001110011100111010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100100111001110011110101101010100101001010011100111001110011100111001110010100101001010011010110101001110011100111010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101101001010010100101001010011010110101101001000010000100001000010000100011010110101101010100101001010010100101000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101101001010010100101001010011010110101101001000010000100001000010000100011010110101101010100101001010010100101000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101101001010010100101001010011010110101101001000010000100001000010000100011010110101101010100101001010010100101000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111101111011110101001010010100101001010010100111101111011110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111101111011110101001010010100101001010010100111101111011110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111101111011110101001010010100101001010010100111101111011110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110110100101001010010100101001010001101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110110100101001010010100101001010001101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111001110011100111001110011100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111001110011100111001110011100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111001110011100111001110011100110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 9_bonus-godmod
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111101111011110111101111011110110011100111001110011100111100111001110011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111101111011110111101111011110110011100111001110011100111100111001110011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001111101111011110111101111011110110011100111001110011100111100111001110011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111011110111101101001010010100101001010001011010110101100100001000010010100101001010010100101001110111101111010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111011110111101101001010010100101001010001011010110101100100001000010010100101001010010100101001110111101111010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100010110101101011001000010000010000100001001010010100101001011010110101100010000100001001011010110010000100001001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100010110101101011001000010000010000100001001010010100101001011010110101100010000100001001011010110010000100001001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100010110101101011001000010000010000100001001010010100101001011010110101100010000100001001011010110010000100001001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100010100101001010010110101110100101001010000110001100011001011010110101100110001100011001010010100101101011010111010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100010100101001010010110101110100101001010000110001100011001011010110101100110001100011001010010100101101011010111010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100010100101001010010110101110100101001010000110001100011001011010110101100110001100011001010010100101101011010111010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100001110011100111010100101000110001100011001010010100101001011010110101110100101001010000111001110101101011010110001000010000100110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100001110011100111010100101000110001100011001010010100101001011010110101110100101001010000111001110101101011010110001000010000100110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100001110011100111010100101000110001100011001010010100101001011010110101110100101001010000111001110101101011010110001000010000100110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100010100101001010010100101010100101001010001010010100101001010010100101010100101001010010001100010101101011010111110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101101001010010100010100101001010010100101010100101001010001010010100101001010010100101010100101001010010001100010101101011010111110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111011110111101101001010010100101001010010100111001110000010000100001000010000100001000110001100011010100101001010010100101001010010100101001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111011110111101101001010010100101001010010100111001110000010000100001000010000100001000110001100011010100101001010010100101001010010100101001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111011110111101101001010010100101001010010100111001110000010000100001000010000100001000110001100011010100101001010010100101001010010100101001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010110101101011000010000100001111011110111101111001110001010010100101001010010100101010001100011000100111001110011110001100011010010100101001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010110101101011000010000100001111011110111101111001110001010010100101001010010100101010001100011000100111001110011110001100011010010100101001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010110101101011000010000100001111011110111101111001110001010010100101001010010100101010001100011000100111001110011110001100011010010100101001110111101111010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010100101001010010110101101011010110101101011111011110100111001110011101010010100101000111001110011101011010110101101011010110101001010010101110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010100101001010010110101101011010110101101011111011110100111001110011101010010100101000111001110011101011010110101101011010110101001010010101110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010100101001010010110101101011010110101101011111011110100111001110011101010010100101000111001110011101011010110101101011010110101001010010101110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111001110011100010100101001010011110111101111010110101101011010110101101110011100111010100101001010001010010100101001011010110101101011010111110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111001110011100010100101001010011110111101111010110101101011010110101101110011100111010100101001010001010010100101001011010110101101011010111110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111001110011100010100101001010011110111101111010110101101011010110101101110011100111010100101001010001010010100101001011010110101101011010111110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100001100011000110010100101001010100101001000001000010000101011010110101110100101001010001010010100101001011010111000110001100011010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100001100011000110010100101001010100101001000001000010000101011010110101110100101001010001010010100101001011010111000110001100011010010100101000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100001100011000110010100101001011010110101101011010110101100010000100001001010010100101001010010100011000110001101110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100001100011000110010100101001011010110101101011010110101100010000100001001010010100101001010010100011000110001101110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100001100011000110010100101001011010110101101011010110101100010000100001001010010100101001010010100011000110001101110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111001110011100001100011001010010100101001011010110101110100101001010001010010100101001010010101110011100111000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111001110011100001100011001010010100101001011010110101110100101001010001010010100101001010010101110011100111000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111001110011100001100011001010010100101001011010110101110100101001010001010010100101001010010101110011100111000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010000111001110011101010010100101000110001100011011110111101111000110001100110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010000111001110011101010010100101000110001100011011110111101111000110001100110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010000111001110011101010010100101000110001100011011110111101111000110001100110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111001110011100111011110101010010100101001010010100101001011010110101101011010110101110001100011110011100111000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101111001110011100111011110101010010100101001010010100101001011010110101101011010110101110001100011110011100111000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011101001010010100111001110000110001100011000010000100001000010000100001000110001100011000110001101010010100101001001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011101001010010100111001110000110001100011000010000100001000010000100001000110001100011000110001101010010100101001001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011101001010010100111001110000110001100011000010000100001000010000100001000110001100011000110001101010010100101001001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 10_bonus-wallhack
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111100111001110011100111001100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111100111001110011100111001100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111100111001110011100111001100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001010000100001000010000100001001000010000100010110101101011010110101101011111001110011100111001110011101111011110111100111001110011100111001110011100111001110011100111001110111101111011110011100111001110011100100111001110011001010010100101"),
                ("0010100101001010000100001000010000100001001000010000100010110101101011010110101101011111001110011100111001110011101111011110111100111001110011100111001110011100111001110011100111001110111101111011110011100111001110011100100111001110011001010010100101"),
                ("0010100101001010000100001000010000100001001000010000100010110101101011010110101101011111001110011100111001110011101111011110111100111001110011100111001110011100111001110011100111001110111101111011110011100111001110011100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110000100001000010011000110000011000110001110111101111011100011000110001110100101001010001100011000001100011000111011110111101110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110000100001000010011000110000011000110001110111101111011100011000110001110100101001010001100011000001100011000111011110111101110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110000100001000010011000110000011000110001110111101111011100011000110001110100101001010001100011000001100011000111011110111101110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110010110101101001000010000100010110101101011100001000010000010110101101011010110101100011000110001100011000110001110100101001010001100011000001100011000110001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110010110101101001000010000100010110101101011100001000010000010110101101011010110101100011000110001100011000110001110100101001010001100011000001100011000110001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110010110101101001000010000100010110101101011100001000010000010110101101011010110101100011000110001100011000110001110100101001010001100011000001100011000110001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110001100011000110011000110001100011000110001100011000110001100011000110010100101001010001100011000110001100011000110001100011000110001100011001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110001100011000110011000110001100011000110001100011000110001100011000110010100101001010001100011000110001100011000110001100011000110001100011001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110010000100001000010000100001010010100101001010010100101100001000000000000000000000000000000000010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110010000100001000010000100001010010100101001010010100101100001000000000000000000000000000000000010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110010000100001000010000100001010010100101001010010100101100001000000000000000000000000000000000010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110001100011000110001100011000010000100001001100011000110000011000110001110111101111011100011000111010010100101000001100011000110010100101001011010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110001100011000110001100011000010000100001001100011000110000011000110001110111101111011100011000111010010100101000001100011000110010100101001011010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110001100011000110001100011000010000100001001100011000110000011000110001110111101111011100011000111010010100101000001100011000110010100101001011010010100110011100111001001010010100101"),
                ("0010100101001010000100001000010010000100001000010000100001010010100101010110101101011010110101101011010110101101011010110101100011000110001100011000110001100011000111010010100101000001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001010000100001000010010000100001000010000100001010010100101010110101101011010110101101011010110101101011010110101100011000110001100011000110001100011000111010010100101000001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001010000100001000010010000100001000010000100001010010100101010110101101011010110101101011010110101101011010110101100011000110001100011000110001100011000111010010100101000001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110011000110001100011000110000010000100001001100011000110001100011000110001100011000110001100011001010010100101000110001100011000110001100011001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110011000110001100011000110000010000100001001100011000110001100011000110001100011000110001100011001010010100101000110001100011000110001100011001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110011000110001100011000110000010000100001001100011000110001100011000110001100011000110001100011001010010100101000110001100011000110001100011001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110010000100001000010000100100001000010000000000000000000000000000010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110010000100001000010000100100001000010000000000000000000000000000010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110011000110001100000110001100011000110001110111101111011100011000110001110100101001010001100011000001100011000111011110111101110001100011000111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110011000110001100000110001100011000110001110111101111011100011000110001110100101001010001100011000001100011000111011110111101110001100011000111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111101111011110011000110001100000110001100011000110001110111101111011100011000110001110100101001010001100011000001100011000111011110111101110001100011000111010010100100111001110011001010010100101"),
                ("0010100101001010000100001000010010000100001000010000100010110101101011010110101101011010110101100011000110001100011000110001100011000110001110100101001010001100011000001100011000110001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001010000100001000010010000100001000010000100010110101101011010110101101011010110101100011000110001100011000110001100011000110001110100101001010001100011000001100011000110001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001010000100001000010010000100001000010000100010110101101011010110101101011010110101100011000110001100011000110001100011000110001110100101001010001100011000001100011000110001100011000110001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111111111111111001100011000110001100011011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111111111111111001100011000110001100011011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111111111111111001100011000110001100011011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100100111001110011001010010100101"),
                ("0010100101001011100111001110010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011100111001110010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 11_bonus-speed
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110110100101001010001100011000110001100011000110001100011000110001100011000110001100011000110001100011001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110110100101001010001100011000110001100011000110001100011000110001100011000110001100011000110001100011001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111100111001110000011000110001100001000010000101011010110101110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111100111001110000011000110001100001000010000101011010110101110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111100111001110000011000110001100001000010000101011010110101110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101111011110101000010000100001000010000100001001010010100111010110101101010000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101111011110101000010000100001000010000100001001010010100111010110101101010000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101111011110101000010000100001000010000100001001010010100111010110101101010000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111101111011110110001100011000110001100011000110001100011000110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111101111011110110001100011000110001100011000110001100011000110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110111101111011110110001100011000110001100011000110001100011000110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101111001110001001010010100101000010000100011000110001100010011100111001110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101111001110001001010010100101000010000100011000110001100010011100111001110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100101001010010100101001010011101111011110110001100011000110001100011000110001100011000110000100000101001010010101110111101111011110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100101001010010100101001010011101111011110110001100011000110001100011000110001100011000110000100000101001010010101110111101111011110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100101001010010100101001010011101111011110110001100011000110001100011000110001100011000110000100000101001010010101110111101111011110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100111011110111101010110101101011000010000100100001000010001011010110101101011010110101101011010110101110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100111011110111101010110101101011000010000100100001000010001011010110101101011010110101101011010110101110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100111011110111101010110101101011000010000100100001000010001011010110101101011010110101101011010110101110000100000101001010010100011000110001101110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110010110101101011000010000100001010110101101011010110101101011010110101101011010110101110000100001000001010010100101001010010100101001010010101111111111111111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110010110101101011000010000100001010110101101011010110101101011010110101101011010110101110000100001000001010010100101001010010100101001010010101111111111111111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110010110101101011000010000100001010110101101011010110101101011010110101101011010110101110000100001000001010010100101001010010100101001010010101111111111111111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010100101001010010110101101011111011110111101101001010010000100001000010000100001000001010010100101001010010100101011101111011010010100101000011000110001101111111111111111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010100101001010010110101101011111011110111101101001010010000100001000010000100001000001010010100101001010010100101011101111011010010100101000011000110001101111111111111111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100010100101001010010110101101011111011110111101101001010010000100001000010000100001000001010010100101001010010100101011101111011010010100101000011000110001101111111111111111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110111011110111101010000100001000010000100011100111001110011101111011110100110001100011011101111011110101000010000100001000010001110011100111001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110111011110111101010000100001000010000100011100111001110011101111011110100110001100011011101111011110101000010000100001000010001110011100111001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100010000100001000011110111101111011100111001000010000100010100101001010010100101001010001000010000100001111011110111001110011100100001000010001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100010000100001000011110111101111011100111001000010000100010100101001010010100101001010001000010000100001111011110111001110011100100001000010001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100010000100001000011110111101111011100111001000010000100010100101001010010100101001010001000010000100001111011110111001110011100100001000010001010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111011110111101010000100001000011100111001110111101111011000110001100010100101001010011100111001110001000010000100001110011101111011110111101100011000110001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111011110111101010000100001000011100111001110111101111011000110001100010100101001010011100111001110001000010000100001110011101111011110111101100011000110001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111011110111101010000100001000011100111001110111101111011000110001100010100101001010011100111001110001000010000100001110011101111011110111101100011000110001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111011110111101010000100001000110001100011100111001110001101011010110101101011010110111101111011110101000010001100011000110001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111011110111101010000100001000110001100011100111001110001101011010110101101011010110111101111011110101000010001100011000110001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111011110111101010000100001000110001100011100111001110001101011010110101101011010110111101111011110101000010001100011000110001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101101001010010100101001010001101011010110101101011010110101101011010110101101011010110110100101001010010100101000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101101001010010100101001010001101011010110101101011010110101101011010110101101011010110110100101001010010100101000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011110011100111001110011100110011100111001110011100111001110011100111001110011100111001111001110011100111001110011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011110011100111001110011100110011100111001110011100111001110011100111001110011100111001111001110011100111001110011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011110011100111001110011100110011100111001110011100111001110011100111001110011100111001111001110011100111001110011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 12_bonus-addbomb
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111100111001110011100111001110011001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111100111001110011100111001110011001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111100111001110011100111001110011001110011100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010011100111001111111111111111110111101111011010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010011100111001111111111111111110111101111011010010100101000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011101111011110111100111001110011100111001110001111011110111111101111010111001110011100010000100001001001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011101111011110111100111001110011100111001110001111011110111111101111010111001110011100010000100001001001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011101111011110111100111001110011100111001110001111011110111111101111010111001110011100010000100001001001110011100111010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000111011110111101011110111101111011110111111100111001110000101001010010100100001000010011101111010010000100001000010100101001011110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000111011110111101011110111101111011110111111100111001110000101001010010100100001000010011101111010010000100001000010100101001011110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000111011110111101011110111101111011110111111100111001110000101001010010100100001000010011101111010010000100001000010100101001011110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100111011110111101010110101101011000010000110000100001000010100101001010000001000010000101011010110101100010000101010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100111011110111101010110101101011000010000110000100001000010100101001010000001000010000101011010110101100010000101010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100111011110111101010110101101011000010000110000100001000010100101001010000001000010000101011010110101100010000101010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111011110111101011110111101111000010000100001001000010010000100001000010100101001010010000100001000010000100001000001111011111110011100111001110011100111001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111011110111101011110111101111000010000100001001000010010000100001000010100101001010010000100001000010000100001000001111011111110011100111001110011100111001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111100001000010000010110101101011100001000001111011110111111101111011110110100101001010001111011110111101110011101110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111100001000010000010110101101011100001000001111011110111111101111011110110100101001010001111011110111101110011101110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111100001000010000010110101101011100001000001111011110111111101111011110110100101001010001111011110111101110011101110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111100001000010000100001000010000011110111101111011110111101111011110111111101111011110110100101001010010100101001010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111100001000010000100001000010000011110111101111011110111101111011110111111101111011110110100101001010010100101001010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111100001000010000100001000010000011110111101111011110111101111011110111111101111011110110100101001010010100101001010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111111101111011110111101111011110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111111101111011110111101111011110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011110111101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111111101111011110111101111011110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110011110111101111011110111101111011110111101111011110111101111011110111101110011100111011101111011110111101111011010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110011110111101111011110111101111011110111101111011110111101111011110111101110011100111011101111011110111101111011010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100001100011000110011110111101111011110111101111011110111101111011110111101111011110111101110011100111011101111011110111101111011010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111001110011100111011110111101011110111101111011110111101111011110111101110011100111011101111011110101110011100111011101111011010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111001110011100111011110111101011110111101111011110111101111011110111101110011100111011101111011110101110011100111011101111011010010100101001010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100101001010010100111011110111101011100111001110011100111011101111011110111101111011110111101111011110110100101001010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100101001010010100111011110111101011100111001110011100111011101111011110111101111011110111101111011110110100101001010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100101001010010100111011110111101011100111001110011100111011101111011110111101111011110111101111011110110100101001010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000101001010010100111011110111101111011110111101111011110110100101001010010100101001010010100101001010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000101001010010100111011110111101111011110111101111011110110100101001010010100101001010010100101001010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000101001010010100111011110111101111011110111101111011110110100101001010010100101001010010100101001010010100101001010010100101001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010010100101000110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010010100101000110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 13_bonus-power
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110101100011000110001101011010110101101011010110101100011000110101101011010110101101011010110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101101011010110101100011000110001101011010110101101011010110101100011000110101101011010110101101011010110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101100011000110011010110101101001100011000110001100011000110001000010000110001100011000110001100011001100011000110000110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101100011000110011010110101101001100011000110001100011000110001000010000110001100011000110001100011001100011000110000110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011010110101100011000110011010110101101001100011000110001100011000110001000010000110001100011000110001100011001100011000110000110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011000110001100011000110001001010010100101000010000100001100011000110001000010000100001000010000110001100011000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011000110001100011000110001001010010100101000010000100001100011000110001000010000100001000010000110001100011000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011000110001100011000110001001010010100101000010000100001100011000110001000010000100001000010000110001100011000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011000110001100110001100011000000010000100001000010000101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011000110001100110001100011000000010000100001000010000101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011000110001100110001100011000000010000100001000010000101000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100110001100011000000010000100001000010000101000010000100001000010000100000001000010000101000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100110001100011000000010000100001000010000101000010000100001000010000100000001000010000101000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100101111011110111010000100001000111011110110111101111011101000010000100011101111011110100100001000010001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100101111011110111010000100001000111011110110111101111011101000010000100011101111011110100100001000010001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100101111011110111010000100001000111011110110111101111011101000010000100011101111011110100100001000010001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010010100101001010000100001000010000100001000101001010000001000010000101000010000100010100101001010000100001000010001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010010100101001010000100001000010000100001000101001010000001000010000101000010000100010100101001010000100001000010001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010010100101001010000100001000010000100001000101001010000001000010000101000010000100010100101001010000100001000010001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000010000100001000111101111000001000010000101000010000100011101111011110100001000010000101000010000100001000010000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000010000100001000111101111000001000010000101000010000100011101111011110100001000010000101000010000100001000010000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000010000100001000111101111000001000010000101000010000100011101111011110100001000010000101000010000100001000010000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000001000010000100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000001000010000100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000001000010000100010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111100111001010010100101001010000100001000011000110001100101001010010100101001010010100101001010010100101001010010100101001010001000010000100001000010000100101001010010110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111100111001010010100101001010000100001000011000110001100101001010010100101001010010100101001010010100101001010010100101001010001000010000100001000010000100101001010010110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100110001100011000010000100001000010000100001000011000110011001110011100111001110011100110100101001010011000110001100001000010000100001000010001101011010110100110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100110001100011000010000100001000010000100001000011000110011001110011100111001110011100110100101001010011000110001100001000010000100001000010001101011010110100110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100110001100011000010000100001000010000100001000011000110011001110011100111001110011100110100101001010011000110001100001000010000100001000010001101011010110100110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100110101101011010010000100001000010000100001100011000110001100011000110001001010010100101000010000100001000010001101011010110100110001100011000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100110101101011010010000100001000010000100001100011000110001100011000110001001010010100101000010000100001000010001101011010110100110001100011000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100110101101011010010000100001000010000100001100011000110001100011000110001001010010100101000010000100001000010001101011010110100110001100011000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011000110001100011000110001100010000100001000010000100001000010000100001000010000100001001010010100101100011000110001100011000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011000110001100011000110001100010000100001000010000100001000010000100001000010000100001001010010100101100011000110001100011000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011000110001100011000110001100010000100001000010000100001000010000100001000010000100001001010010100101100011000110001100011000110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011000110001100011000110001100011000110001100011000110001100011000110001101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101011000110001100011000110001100011000110001100011000110001100011000110001101011010110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 14_malus-inversed-commands
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010110011100111001110011100111001110011100111001110011100111001110011100111001101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111110011100111001110011100111001110011100111001110011100111001110011100111001100101"),
                ("0010110011100111001110011100111001110011100111001110011100111001110011100111001101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111110011100111001110011100111001110011100111001110011100111001110011100111001100101"),
                ("0010110011100111001110011100111001110011100111001110011100111001110011100111001101111011110111101111011110111101111011110111101111011110111101111011110111101111011110111110011100111001110011100111001110011100111001110011100111001110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101101011010110110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101011010110101101111011110111110011100111001100101"),
                ("0010101111011110111101011010110101101111011110111101111011110111101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101111011110111101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101111011110111101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101111011110111101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101111011110111101111011110111101111011110111101011010110101101011010110101101011010110101101011010110101101111011110111101111011110111101111011110111101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101011010110101101111011110111101111011110111101111011110111101011010110101101011010110101101111011110111101111011110111101111011110111101011010110101101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101011010110101101111011110111101111011110111101111011110111101011010110101101011010110101101111011110111101111011110111101111011110111101011010110101101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101011010110101101111011110111101111011110111101111011110111101011010110101101011010110101101111011110111101111011110111101111011110111101011010110101101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101111011110111101111011110111110100101001010001111011110111110100101001010010100101001010001111011110111110100101001010001111011110111101111011110111101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101111011110111101111011110111110100101001010001111011110111110100101001010010100101001010001111011110111110100101001010001111011110111101111011110111101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101111011110111101111011110111101111011110111110100101001010001111011110111110100101001010010100101001010001111011110111110100101001010001111011110111101111011110111101111011110111101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101011010110101101111011110111101111011110111110100101001010001011010110101110100101001010010100101001010001011010110101110100101001010001111011110111101111011110111101011010110101101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101011010110101101111011110111101111011110111110100101001010001011010110101110100101001010010100101001010001011010110101110100101001010001111011110111101111011110111101011010110101101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101011010110101101111011110111101111011110111110100101001010001011010110101110100101001010010100101001010001011010110101110100101001010001111011110111101111011110111101011010110101101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101011010110101101011010110101101011010110101110100101001010010100101001010010100101001010010100101001010010100101001010010100101001010001011010110101101011010110101101011010110101101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101011010110101101011010110101101011010110101110100101001010010100101001010010100101001010010100101001010010100101001010010100101001010001011010110101101011010110101101011010110101101011010110101101111011110111100101"),
                ("0010101111011110111101011010110101101011010110101101011010110101101011010110101110100101001010010100101001010010100101001010010100101001010010100101001010010100101001010001011010110101101011010110101101011010110101101011010110101101111011110111100101"),
                ("0010110011100111001101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101110100101001010010100101001010001011010110101101011010110101101011010110101101011010110101101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101110100101001010010100101001010001011010110101101011010110101101011010110101101011010110101101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101111011110111101011010110101101011010110101101011010110101101011010110101101011010110101110100101001010010100101001010001011010110101101011010110101101011010110101101011010110101101011010110101101111011110111110011100111001100101"),
                ("0010110011100111001101101011010110101111011110111101111011110111101011010110101101011010110101101011010110101110100101001010010100101001010001011010110101101011010110101101011010110101101111011110111101111011110111101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101111011110111101111011110111101011010110101101011010110101101011010110101110100101001010010100101001010001011010110101101011010110101101011010110101101111011110111101111011110111101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101111011110111101111011110111101011010110101101011010110101101011010110101110100101001010010100101001010001011010110101101011010110101101011010110101101111011110111101111011110111101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101011010110101110100101001010010100101001010010100101001010010100101001010010100101001010010100101001010001011010110101101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101011010110101110100101001010010100101001010010100101001010010100101001010010100101001010010100101001010001011010110101101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101011010110101110100101001010010100101001010010100101001010010100101001010010100101001010010100101001010001011010110101101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101011010110101110100101001010001011010110101101111011110111101111011110111101011010110101110100101001010001011010110101101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101011010110101110100101001010001011010110101101111011110111101111011110111101011010110101110100101001010001011010110101101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111101011010110101110100101001010001011010110101101111011110111101111011110111101011010110101110100101001010001011010110101101111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111110100101001010010100101001010001111011110111101111011110111101111011110111101111011110111110100101001010010100101001010001111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111110100101001010010100101001010001111011110111101111011110111101111011110111101111011110111110100101001010010100101001010001111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001101101011010110101101011010110101111011110111110100101001010010100101001010001111011110111101111011110111101111011110111101111011110111110100101001010010100101001010001111011110111101101011010110101101011010110110011100111001100101"),
                ("0010110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001100101"),
                ("0010110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001100101"),
                ("0010110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 15_malus-disable-bombs
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011110011100111001110011100111001100111001110011100111001111001110011100110100101001010010100101001010011001110011100110011100111001110011100111100111001110011100111001110011001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011110011100111001110011100111001100111001110011100111001111001110011100110100101001010010100101001010011001110011100110011100111001110011100111100111001110011100111001110011001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011110011100111001110011100111001100111001110011100111001111001110011100110100101001010010100101001010011001110011100110011100111001110011100111100111001110011100111001110011001110011100111001110011001010010100101"),
                ("0010100101001011100111001110011010010100101001010010100101001010010100111011110111101101001010010100101001010001000010000100000011000110001110100101001010010100101001110111101111011010010100101001010010100101001010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100101001010010100101001010010100111011110111101101001010010100101001010001000010000100000011000110001110100101001010010100101001110111101111011010010100101001010010100101001010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010000100001000000110001100011111001110011100001110011100111001110011100001000010000101000010000100011101111011110100000000001010010100101000001100011000110100001000010001010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010000100001000000110001100011111001110011100001110011100111001110011100001000010000101000010000100011101111011110100000000001010010100101000001100011000110100001000010001010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010000100001000000110001100011111001110011100001110011100111001110011100001000010000101000010000100011101111011110100000000001010010100101000001100011000110100001000010001010010100110011100111001001010010100101"),
                ("0010100101001011001110011100111010010100000110001100011001110011100111100001000010000111011110100011000110001100001000010000101000010000100000011000110001110100101000000000000000001110111101111010001100011000111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100000110001100011001110011100111100001000010000111011110100011000110001100001000010000101000010000100000011000110001110100101000000000000000001110111101111010001100011000111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100000110001100011001110011100111100001000010000111011110100011000110001100001000010000101000010000100000011000110001110100101000000000000000001110111101111010001100011000111010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111110011100111001110011100010110101101011010110101101011101001010000011000110001101000010000100001000010000100000011000110001110100101001110111101111011010010100101001110011100111001110111101100111001110011001010010100101"),
                ("0010100101001011001110011100111110011100111001110011100010110101101011010110101101011101001010000011000110001101000010000100001000010000100000011000110001110100101001110111101111011010010100101001110011100111001110111101100111001110011001010010100101"),
                ("0010100101001011001110011100111110011100111001110011100010110101101011010110101101011101001010000011000110001101000010000100001000010000100000011000110001110100101001110111101111011010010100101001110011100111001110111101100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111111111111111010110101101011000010000100001100001000000011000110001101000010000100001000010000100000011000110001110100101001110111101111011010010100101000000000000000001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100111111111111111010110101101011000010000100001100001000000011000110001101000010000100001000010000100000011000110001110100101001110111101111011010010100101000000000000000001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100100001000010000010110101101011000010000100001000010000101111011110111110100101001010010100101001010011110111101111001110011101110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100100001000010000010110101101011000010000100001000010000101111011110111110100101001010010100101001010011110111101111001110011101110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100100001000010000010110101101011000010000100001000010000101111011110111110100101001010010100101001010011110111101111001110011101110111101111011010010100101001110011100111001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100100001000010000011110111101111011110111101111010110101101011010110101110000100001000010000100001000001111011110111111101111011110011100111001010010100101000000000000000001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100100001000010000011110111101111011110111101111010110101101011010110101110000100001000010000100001000001111011110111111101111011110011100111001010010100101000000000000000001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100100001000010000011110111101111011110111101111010110101101011010110101110000100001000010000100001000001111011110111111101111011110011100111001010010100101000000000000000001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011100111001110000110001100011101001010010100011110111110000100001000010000100001000001111011110111101110011100111010100101001010010100101000001100011000111010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011100111001110000110001100011101001010010100011110111110000100001000010000100001000001111011110111101110011100111010100101001010010100101000001100011000111010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011001110011100111010010100011100111001110000110001100011101001010010100011110111110000100001000010000100001000001111011110111101110011100111010100101001010010100101000001100011000111010010100101001010010100100111001110011001010010100101"),
                ("0010100101001011100111001110011010010100000110001100011000010000100001010000100001000101001010001111011110111101111011110111101110011100111011100111001110010100101000100001000010000000100001000010001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100000110001100011000010000100001010000100001000101001010001111011110111101111011110111101110011100111011100111001110010100101000100001000010000000100001000010001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100000110001100011000010000100001010000100001000101001010001111011110111101111011110111101110011100111011100111001110010100101000100001000010000000100001000010001100011000111010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100000010000100001000010000100001010000100001000101001010011101111011110111101111011110111101111011110110100101001010010100101000100001000010000000100001000010000100001000011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100000010000100001000010000100001010000100001000101001010011101111011110111101111011110111101111011110110100101001010010100101000100001000010000000100001000010000100001000011010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010000100001000000110001100011000110001100011101001010010100101001010010100101001010010100101001010010100101001010010100101000001100011000110001100011000110100001000010001010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010000100001000000110001100011000110001100011101001010010100101001010010100101001010010100101001010010100101001010010100101000001100011000110001100011000110100001000010001010010100110011100111001001010010100101"),
                ("0010100101001011100111001110011010010100010000100001000000110001100011000110001100011101001010010100101001010010100101001010010100101001010010100101001010010100101000001100011000110001100011000110100001000010001010010100110011100111001001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101000000000000000001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101000000000000000001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101111001110011100000000000000000101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101000000000000000001110011100111000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111000110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010010100101000110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011010110101101011010110101101011010110101101101001010010100101001010010100101001010010100101001010010100101001010010100101000110101101011010110101101011010110101101011010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),

                -- 16_malus-remove-power
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011011010110101101011010110101101011010110101101011010110101100011000110001101011010110101101011010110101100011000110001100011001001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011011010110101101011010110101101011010110101101011010110101100011000110001101011010110101101011010110101100011000110001100011001001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011011010110101101011010110101100011000110011010110101101001100011000110001100011000110011000110001001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011011010110101101011010110101100011000110011010110101101001100011000110001100011000110011000110001001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011011010110101101011010110101100011000110011010110101101001100011000110001100011000110011000110001001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011011000110001001010010100101000010000100001100011000110001001010010100110011100111001110011100111001110011100111001110011100111100111001100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011011000110001001010010100101000010000100001100011000110001001010010100110011100111001110011100111001110011100111001110011100111100111001100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011011000110001001010010100101000010000100001100011000110001001010010100110011100111001110011100111001110011100111001110011100111100111001100111001110011001010010100101"),
                ("0010100101001011001110011100111111011110100111001110011100111001110011100111001110011100111001110111101111011101000010000100001001010010100110011100111001110011100111001110011100111001110011100110100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111111011110100111001110011100111001110011100111001110011100111001110111101111011101000010000100001001010010100110011100111001110011100111001110011100111001110011100110100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111111011110100111001110011100111001110011100111001110011100111001110111101111011101000010000100001001010010100110011100111001110011100111001110011100111001110011100110100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101110011100111001100111001110011100111001110011100111001110011100111001101001010010100110011100111001110011100111001110011100111001110011100110100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101110011100111001100111001110011100111001110011100111001110011100111001101001010010100110011100111001110011100111001110011100111001110011100110100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100101011010110101100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100101011010110101100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110101101011000110001100101011010110101100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010010100101001010000100001000010010100101001100111001110011100111001110011100111001110011100111001110011100111001101000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010010100101001010000100001000010010100101001100111001110011100111001110011100111001110011100111001110011100111001101000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010010100101001010000100001000010010100101001100111001110011100111001110011100111001110011100111001110011100111001101000010000100001000010000100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000010000100001000100111001110011100111001110011100111001110011100111001110011100111001101001010010100001000010000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000010000100001000100111001110011100111001110011100111001110011100111001110011100111001101001010010100001000010000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000010000100001000100111001110011100111001110011100111001110011100111001110011100111001101001010010100001000010000100001000010000100101001010011100111001100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110100101001010010100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110100101001010010100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100010000100001000010000100001000100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100110100101001010010100001000010000100101001010010110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111100111001010010100101001100111001110011100111001110011100111001110011100111001101100011000110010011100111001110011100111001110011100111001110011100111101011010110100110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111100111001010010100101001100111001110011100111001110011100111001110011100111001101100011000110010011100111001110011100111001110011100111001110011100111101011010110100110001100011000110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100100111001110011100111001110011100111001110011100111001110011100111001111001110011100110100101001010010011100111001110011100111001110011100111001110011100111100111001110010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100100111001110011100111001110011100111001110011100111001110011100111001111001110011100110100101001010010011100111001110011100111001110011100111001110011100111100111001110010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100110110001100100111001110011100111001110011100111001110011100111001110011100111001111001110011100110100101001010010011100111001110011100111001110011100111001110011100111100111001110010110101101100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011010010100101100011000110001100011000110001001010010100101000010000100010011100111001110011100111001110011100111001110011100110110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011010010100101100011000110001100011000110001001010010100101000010000100010011100111001110011100111001110011100111001110011100110110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011010010100101100011000110001100011000110001001010010100101000010000100010011100111001110011100111001110011100111001110011100110110001100100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011110011100111001010000100001000010000100001000010000100001000010000100001001010010100101100011001001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011110011100111001010000100001000010000100001000010000100001000010000100001001010010100101100011001001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011110011100111001010000100001000010000100001000010000100001000010000100001001010010100101100011001001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011011000110001100011010110101101011000110001100011000110001100011000110001100011000110001100011000110001101011010110101101011011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011011000110001100011010110101101011000110001100011000110001100011000110001100011000110001100011000110001101011010110101101011011001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001011001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011100111001110011001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101"),
                ("0010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101001010010100101")
            );
    end init_mem;

    constant rom : memory_t := init_mem;
    signal real_row : integer range 0 to 2051 := 0;
    signal out_color_reg : std_logic_vector(49 downto 0) := (others => '0');
begin
    process(in_sprite_id, in_sprite_row, in_sprite_col)
    begin
        case in_sprite_id is
            when 1 => real_row <= in_sprite_row;
            when 2 => real_row <= 50 + in_sprite_row;
            when 3 => real_row <= 100 + in_sprite_row;
            when 4 =>
                case in_sprite_state is
                    when 0 => real_row <= 150 + in_sprite_row;
                    when others => null;
                end case;
            when 5 =>
                case in_sprite_state is
                    when 0 => real_row <= 202 + in_sprite_row;
                    when 1 => real_row <= 252 + in_sprite_row;
                    when 2 => real_row <= 302 + in_sprite_row;
                    when 3 => real_row <= 352 + in_sprite_row;
                    when others => null;
                end case;
            when 6 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 402 + in_sprite_row;
                            when D_LEFT => real_row <= 452 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 502 + in_sprite_row;
                            when D_LEFT => real_row <= 552 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 602 + in_sprite_row;
                            when D_LEFT => real_row <= 652 + in_sprite_row;
                            when others => null;
                        end case;
                    when 3 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 702 + in_sprite_row;
                            when D_LEFT => real_row <= 752 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 7 =>
                case in_sprite_state is
                    when 0 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 802 + in_sprite_row;
                            when D_LEFT => real_row <= 852 + in_sprite_row;
                            when D_DOWN => real_row <= 902 + in_sprite_row;
                            when D_RIGHT => real_row <= 952 + in_sprite_row;
                            when others => null;
                        end case;
                    when 1 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1002 + in_sprite_row;
                            when D_LEFT => real_row <= 1052 + in_sprite_row;
                            when D_DOWN => real_row <= 1102 + in_sprite_row;
                            when D_RIGHT => real_row <= 1152 + in_sprite_row;
                            when others => null;
                        end case;
                    when 2 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1202 + in_sprite_row;
                            when D_LEFT => real_row <= 1252 + in_sprite_row;
                            when D_DOWN => real_row <= 1302 + in_sprite_row;
                            when D_RIGHT => real_row <= 1352 + in_sprite_row;
                            when others => null;
                        end case;
                    when 3 =>
                        case in_sprite_direction is
                            when D_UP => real_row <= 1402 + in_sprite_row;
                            when D_LEFT => real_row <= 1452 + in_sprite_row;
                            when D_DOWN => real_row <= 1502 + in_sprite_row;
                            when D_RIGHT => real_row <= 1552 + in_sprite_row;
                            when others => null;
                        end case;
                    when others => null;
                end case;
            when 8 => real_row <= 1602 + in_sprite_row;
            when 9 => real_row <= 1652 + in_sprite_row;
            when 10 => real_row <= 1702 + in_sprite_row;
            when 11 => real_row <= 1752 + in_sprite_row;
            when 12 => real_row <= 1802 + in_sprite_row;
            when 13 => real_row <= 1852 + in_sprite_row;
            when 14 => real_row <= 1902 + in_sprite_row;
            when 15 => real_row <= 1952 + in_sprite_row;
            when 16 => real_row <= 2002 + in_sprite_row;
            when others => null;
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            out_color_reg <= rom(real_row);
        end if;
    end process;
    out_color <= out_color_reg(((in_sprite_col + 1) * 5 - 1) downto (in_sprite_col * 5));
end behavioural;
